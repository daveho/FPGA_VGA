// Testbench for vcount module

`include "testbench.vh"

module vcount_tb();

  `include "timing.vh"

  integer k;

  // helper task to generate a specified number of clock pulses
  task automatic genclock( input [11:0] ticks, output clk ); begin
    for ( k = 0; k < ticks; k++ ) begin
      clk = 1;
      #1;
      clk = 0;
      #1;
    end
  end endtask

  // The testbench just needs to control -RST and CLK
  reg nrst, clk;

  // Outputs generated by the hcount module
  wire hCountEnd, hBeginPulse, hEndPulse, hVisEnd, hBeginActive, hEndActive;

  // Outputs generated by the vcount module
  wire vCountZero, vBeginPulse, vEndPulse, vVisEnd, vCountEnd, vEndActive;
  wire [11:0] vCount;

  // Instantiate hcount module
  hcount hcount_instance( // Inputs
                          .nrst( nrst ),
                          .clk( clk ),
                          // Outputs
                          .hCountEnd( hCountEnd ),
                          .hBeginPulse( hBeginPulse ),
                          .hEndPulse( hEndPulse ),
                          .hVisEnd( hVisEnd ),
                          .hBeginActive( hBeginActive ),
                          .hEndActive( hEndActive ) );

  // Instantiate vcount module. Note that the hEndPulse signal
  // is used to generate the vCountIncr input to the vcount
  // module.
  vcount vcount_instance( // Inputs
                          .nrst( nrst ),
                          .clk( clk ),
                          .vCountIncr( hEndPulse ),
                          .hCountEnd( hCountEnd ),
                          // Outputs
                         .vCountZero( vCountZero ),
                         .vBeginPulse( vBeginPulse ),
                         .vEndPulse( vEndPulse ),
                         .vVisEnd( vVisEnd ),
                         .vCountEnd( vCountEnd ),
                         .vEndActive( vEndActive ),
                         .vCount( vCount ) );

  initial begin
    // generate dump file we can inspect using gtkwave
    $dumpfile( "vcount_tb.vcd" );
    $dumpvars;
  end

  integer i; // loop counter

  initial begin
    // generate a reset pulse
    nrst = 0;
    clk = 0;
    #1;
    clk = 1;
    #1;
    nrst = 1;
    clk = 0;
    #1;

    // both hcount and vcount are now out of reset

    $display( "vCount=%d", vCount );
    `ASSERT( vCount == V_COUNT_INITIAL_VAL );

    // generate enough ticks to take us to the end of the hsync pulse:
    // this is just before the vertical count will be incremented
    genclock( H_END_PULSE, clk );
    $display( "vCount=%d", vCount );
    `ASSERT( vCount == V_COUNT_INITIAL_VAL );

    // generate one clock pulse: this should increment the vertical count
    genclock( 1, clk );
    $display( "vCount=%d", vCount );
    `ASSERT( vCount == V_COUNT_INITIAL_VAL + 12'd1 );

  end

endmodule;
