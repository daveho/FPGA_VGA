vramData[13'd0] = 8'd31;
vramData[13'd1] = 8'd199;
vramData[13'd2] = 8'd202;
vramData[13'd3] = 8'd87;
vramData[13'd4] = 8'd252;
vramData[13'd5] = 8'd87;
vramData[13'd6] = 8'd200;
vramData[13'd7] = 8'd151;
vramData[13'd8] = 8'd220;
vramData[13'd9] = 8'd121;
vramData[13'd10] = 8'd220;
vramData[13'd11] = 8'd121;
vramData[13'd12] = 8'd183;
vramData[13'd13] = 8'd121;
vramData[13'd14] = 8'd214;
vramData[13'd15] = 8'd121;
vramData[13'd16] = 8'd223;
vramData[13'd17] = 8'd151;
vramData[13'd18] = 8'd223;
vramData[13'd19] = 8'd151;
vramData[13'd20] = 8'd188;
vramData[13'd21] = 8'd151;
vramData[13'd22] = 8'd214;
vramData[13'd23] = 8'd247;
vramData[13'd24] = 8'd202;
vramData[13'd25] = 8'd247;
vramData[13'd26] = 8'd210;
vramData[13'd27] = 8'd151;
vramData[13'd28] = 8'd202;
vramData[13'd29] = 8'd247;
vramData[13'd30] = 8'd210;
vramData[13'd31] = 8'd247;
vramData[13'd32] = 8'd200;
vramData[13'd33] = 8'd135;
vramData[13'd34] = 8'd164;
vramData[13'd35] = 8'd120;
vramData[13'd36] = 8'd210;
vramData[13'd37] = 8'd135;
vramData[13'd38] = 8'd210;
vramData[13'd39] = 8'd135;
vramData[13'd40] = 8'd210;
vramData[13'd41] = 8'd135;
vramData[13'd42] = 8'd16;
vramData[13'd43] = 8'd135;
vramData[13'd44] = 8'd16;
vramData[13'd45] = 8'd120;
vramData[13'd46] = 8'd230;
vramData[13'd47] = 8'd135;
vramData[13'd48] = 8'd30;
vramData[13'd49] = 8'd135;
vramData[13'd50] = 8'd209;
vramData[13'd51] = 8'd135;
vramData[13'd52] = 8'd16;
vramData[13'd53] = 8'd120;
vramData[13'd54] = 8'd210;
vramData[13'd55] = 8'd120;
vramData[13'd56] = 8'd228;
vramData[13'd57] = 8'd120;
vramData[13'd58] = 8'd30;
vramData[13'd59] = 8'd120;
vramData[13'd60] = 8'd210;
vramData[13'd61] = 8'd120;
vramData[13'd62] = 8'd16;
vramData[13'd63] = 8'd135;
vramData[13'd64] = 8'd16;
vramData[13'd65] = 8'd135;
vramData[13'd66] = 8'd16;
vramData[13'd67] = 8'd247;
vramData[13'd68] = 8'd135;
vramData[13'd69] = 8'd120;
vramData[13'd70] = 8'd248;
vramData[13'd71] = 8'd136;
vramData[13'd72] = 8'd0;
vramData[13'd73] = 8'd88;
vramData[13'd74] = 8'd231;
vramData[13'd75] = 8'd136;
vramData[13'd76] = 8'd0;
vramData[13'd77] = 8'd104;
vramData[13'd78] = 8'd17;
vramData[13'd79] = 8'd136;
vramData[13'd80] = 8'd94;
vramData[13'd81] = 8'd200;
vramData[13'd82] = 8'd94;
vramData[13'd83] = 8'd120;
vramData[13'd84] = 8'd252;
vramData[13'd85] = 8'd120;
vramData[13'd86] = 8'd252;
vramData[13'd87] = 8'd120;
vramData[13'd88] = 8'd252;
vramData[13'd89] = 8'd120;
vramData[13'd90] = 8'd252;
vramData[13'd91] = 8'd120;
vramData[13'd92] = 8'd202;
vramData[13'd93] = 8'd120;
vramData[13'd94] = 8'd202;
vramData[13'd95] = 8'd120;
vramData[13'd96] = 8'd202;
vramData[13'd97] = 8'd120;
vramData[13'd98] = 8'd202;
vramData[13'd99] = 8'd120;
vramData[13'd100] = 8'd202;
vramData[13'd101] = 8'd120;
vramData[13'd102] = 8'd31;
vramData[13'd103] = 8'd120;
vramData[13'd104] = 8'd31;
vramData[13'd105] = 8'd120;
vramData[13'd106] = 8'd31;
vramData[13'd107] = 8'd120;
vramData[13'd108] = 8'd31;
vramData[13'd109] = 8'd120;
vramData[13'd110] = 8'd30;
vramData[13'd111] = 8'd120;
vramData[13'd112] = 8'd16;
vramData[13'd113] = 8'd120;
vramData[13'd114] = 8'd16;
vramData[13'd115] = 8'd168;
vramData[13'd116] = 8'd30;
vramData[13'd117] = 8'd168;
vramData[13'd118] = 8'd30;
vramData[13'd119] = 8'd200;
vramData[13'd120] = 8'd214;
vramData[13'd121] = 8'd120;
vramData[13'd122] = 8'd30;
vramData[13'd123] = 8'd120;
vramData[13'd124] = 8'd248;
vramData[13'd125] = 8'd120;
vramData[13'd126] = 8'd193;
vramData[13'd127] = 8'd136;
vramData[13'd128] = 8'd95;
vramData[13'd129] = 8'd152;
vramData[13'd130] = 8'd213;
vramData[13'd131] = 8'd120;
vramData[13'd132] = 8'd197;
vramData[13'd133] = 8'd120;
vramData[13'd134] = 8'd210;
vramData[13'd135] = 8'd120;
vramData[13'd136] = 8'd198;
vramData[13'd137] = 8'd120;
vramData[13'd138] = 8'd164;
vramData[13'd139] = 8'd135;
vramData[13'd140] = 8'd30;
vramData[13'd141] = 8'd135;
vramData[13'd142] = 8'd80;
vramData[13'd143] = 8'd135;
vramData[13'd144] = 8'd150;
vramData[13'd145] = 8'd87;
vramData[13'd146] = 8'd16;
vramData[13'd147] = 8'd135;
vramData[13'd148] = 8'd16;
vramData[13'd149] = 8'd87;
vramData[13'd150] = 8'd126;
vramData[13'd151] = 8'd119;
vramData[13'd152] = 8'd219;
vramData[13'd153] = 8'd126;
vramData[13'd154] = 8'd198;
vramData[13'd155] = 8'd55;
vramData[13'd156] = 8'd16;
vramData[13'd157] = 8'd120;
vramData[13'd158] = 8'd213;
vramData[13'd159] = 8'd120;
vramData[13'd160] = 8'd31;
vramData[13'd161] = 8'd247;
vramData[13'd162] = 8'd31;
vramData[13'd163] = 8'd247;
vramData[13'd164] = 8'd36;
vramData[13'd165] = 8'd119;
vramData[13'd166] = 8'd31;
vramData[13'd167] = 8'd87;
vramData[13'd168] = 8'd24;
vramData[13'd169] = 8'd119;
vramData[13'd170] = 8'd196;
vramData[13'd171] = 8'd247;
vramData[13'd172] = 8'd200;
vramData[13'd173] = 8'd247;
vramData[13'd174] = 8'd202;
vramData[13'd175] = 8'd247;
vramData[13'd176] = 8'd202;
vramData[13'd177] = 8'd247;
vramData[13'd178] = 8'd202;
vramData[13'd179] = 8'd247;
vramData[13'd180] = 8'd202;
vramData[13'd181] = 8'd247;
vramData[13'd182] = 8'd70;
vramData[13'd183] = 8'd247;
vramData[13'd184] = 8'd202;
vramData[13'd185] = 8'd151;
vramData[13'd186] = 8'd212;
vramData[13'd187] = 8'd247;
vramData[13'd188] = 8'd202;
vramData[13'd189] = 8'd247;
vramData[13'd190] = 8'd202;
vramData[13'd191] = 8'd247;
vramData[13'd192] = 8'd16;
vramData[13'd193] = 8'd247;
vramData[13'd194] = 8'd200;
vramData[13'd195] = 8'd87;
vramData[13'd196] = 8'd200;
vramData[13'd197] = 8'd135;
vramData[13'd198] = 8'd202;
vramData[13'd199] = 8'd135;
vramData[13'd200] = 8'd210;
vramData[13'd201] = 8'd152;
vramData[13'd202] = 8'd80;
vramData[13'd203] = 8'd135;
vramData[13'd204] = 8'd202;
vramData[13'd205] = 8'd135;
vramData[13'd206] = 8'd164;
vramData[13'd207] = 8'd120;
vramData[13'd208] = 8'd202;
vramData[13'd209] = 8'd120;
vramData[13'd210] = 8'd181;
vramData[13'd211] = 8'd120;
vramData[13'd212] = 8'd210;
vramData[13'd213] = 8'd120;
vramData[13'd214] = 8'd135;
vramData[13'd215] = 8'd120;
vramData[13'd216] = 8'd145;
vramData[13'd217] = 8'd120;
vramData[13'd218] = 8'd210;
vramData[13'd219] = 8'd120;
vramData[13'd220] = 8'd16;
vramData[13'd221] = 8'd135;
vramData[13'd222] = 8'd85;
vramData[13'd223] = 8'd135;
vramData[13'd224] = 8'd67;
vramData[13'd225] = 8'd87;
vramData[13'd226] = 8'd172;
vramData[13'd227] = 8'd135;
vramData[13'd228] = 8'd31;
vramData[13'd229] = 8'd247;
vramData[13'd230] = 8'd200;
vramData[13'd231] = 8'd135;
vramData[13'd232] = 8'd95;
vramData[13'd233] = 8'd120;
vramData[13'd234] = 8'd214;
vramData[13'd235] = 8'd120;
vramData[13'd236] = 8'd95;
vramData[13'd237] = 8'd120;
vramData[13'd238] = 8'd95;
vramData[13'd239] = 8'd120;
vramData[13'd240] = 8'd95;
vramData[13'd241] = 8'd152;
vramData[13'd242] = 8'd240;
vramData[13'd243] = 8'd136;
vramData[13'd244] = 8'd160;
vramData[13'd245] = 8'd136;
vramData[13'd246] = 8'd175;
vramData[13'd247] = 8'd136;
vramData[13'd248] = 8'd171;
vramData[13'd249] = 8'd136;
vramData[13'd250] = 8'd219;
vramData[13'd251] = 8'd131;
vramData[13'd252] = 8'd255;
vramData[13'd253] = 8'd200;
vramData[13'd254] = 8'd32;
vramData[13'd255] = 8'd72;
vramData[13'd256] = 8'd81;
vramData[13'd257] = 8'd136;
vramData[13'd258] = 8'd149;
vramData[13'd259] = 8'd136;
vramData[13'd260] = 8'd240;
vramData[13'd261] = 8'd136;
vramData[13'd262] = 8'd44;
vramData[13'd263] = 8'd120;
vramData[13'd264] = 8'd140;
vramData[13'd265] = 8'd136;
vramData[13'd266] = 8'd219;
vramData[13'd267] = 8'd128;
vramData[13'd268] = 8'd126;
vramData[13'd269] = 8'd136;
vramData[13'd270] = 8'd0;
vramData[13'd271] = 8'd8;
vramData[13'd272] = 8'd255;
vramData[13'd273] = 8'd232;
vramData[13'd274] = 8'd32;
vramData[13'd275] = 8'd200;
vramData[13'd276] = 8'd214;
vramData[13'd277] = 8'd120;
vramData[13'd278] = 8'd210;
vramData[13'd279] = 8'd120;
vramData[13'd280] = 8'd70;
vramData[13'd281] = 8'd120;
vramData[13'd282] = 8'd253;
vramData[13'd283] = 8'd152;
vramData[13'd284] = 8'd96;
vramData[13'd285] = 8'd152;
vramData[13'd286] = 8'd195;
vramData[13'd287] = 8'd152;
vramData[13'd288] = 8'd30;
vramData[13'd289] = 8'd120;
vramData[13'd290] = 8'd16;
vramData[13'd291] = 8'd120;
vramData[13'd292] = 8'd30;
vramData[13'd293] = 8'd120;
vramData[13'd294] = 8'd17;
vramData[13'd295] = 8'd120;
vramData[13'd296] = 8'd210;
vramData[13'd297] = 8'd120;
vramData[13'd298] = 8'd166;
vramData[13'd299] = 8'd135;
vramData[13'd300] = 8'd253;
vramData[13'd301] = 8'd103;
vramData[13'd302] = 8'd39;
vramData[13'd303] = 8'd135;
vramData[13'd304] = 8'd95;
vramData[13'd305] = 8'd247;
vramData[13'd306] = 8'd126;
vramData[13'd307] = 8'd87;
vramData[13'd308] = 8'd248;
vramData[13'd309] = 8'd55;
vramData[13'd310] = 8'd35;
vramData[13'd311] = 8'd119;
vramData[13'd312] = 8'd67;
vramData[13'd313] = 8'd119;
vramData[13'd314] = 8'd198;
vramData[13'd315] = 8'd55;
vramData[13'd316] = 8'd80;
vramData[13'd317] = 8'd120;
vramData[13'd318] = 8'd16;
vramData[13'd319] = 8'd135;
vramData[13'd320] = 8'd210;
vramData[13'd321] = 8'd183;
vramData[13'd322] = 8'd210;
vramData[13'd323] = 8'd183;
vramData[13'd324] = 8'd210;
vramData[13'd325] = 8'd183;
vramData[13'd326] = 8'd210;
vramData[13'd327] = 8'd183;
vramData[13'd328] = 8'd210;
vramData[13'd329] = 8'd183;
vramData[13'd330] = 8'd210;
vramData[13'd331] = 8'd183;
vramData[13'd332] = 8'd16;
vramData[13'd333] = 8'd151;
vramData[13'd334] = 8'd16;
vramData[13'd335] = 8'd55;
vramData[13'd336] = 8'd202;
vramData[13'd337] = 8'd103;
vramData[13'd338] = 8'd202;
vramData[13'd339] = 8'd103;
vramData[13'd340] = 8'd202;
vramData[13'd341] = 8'd103;
vramData[13'd342] = 8'd202;
vramData[13'd343] = 8'd103;
vramData[13'd344] = 8'd202;
vramData[13'd345] = 8'd231;
vramData[13'd346] = 8'd202;
vramData[13'd347] = 8'd231;
vramData[13'd348] = 8'd80;
vramData[13'd349] = 8'd231;
vramData[13'd350] = 8'd214;
vramData[13'd351] = 8'd183;
vramData[13'd352] = 8'd202;
vramData[13'd353] = 8'd151;
vramData[13'd354] = 8'd209;
vramData[13'd355] = 8'd151;
vramData[13'd356] = 8'd210;
vramData[13'd357] = 8'd183;
vramData[13'd358] = 8'd16;
vramData[13'd359] = 8'd183;
vramData[13'd360] = 8'd202;
vramData[13'd361] = 8'd183;
vramData[13'd362] = 8'd202;
vramData[13'd363] = 8'd55;
vramData[13'd364] = 8'd200;
vramData[13'd365] = 8'd135;
vramData[13'd366] = 8'd209;
vramData[13'd367] = 8'd120;
vramData[13'd368] = 8'd202;
vramData[13'd369] = 8'd135;
vramData[13'd370] = 8'd202;
vramData[13'd371] = 8'd135;
vramData[13'd372] = 8'd16;
vramData[13'd373] = 8'd135;
vramData[13'd374] = 8'd202;
vramData[13'd375] = 8'd135;
vramData[13'd376] = 8'd188;
vramData[13'd377] = 8'd135;
vramData[13'd378] = 8'd248;
vramData[13'd379] = 8'd135;
vramData[13'd380] = 8'd248;
vramData[13'd381] = 8'd135;
vramData[13'd382] = 8'd0;
vramData[13'd383] = 8'd151;
vramData[13'd384] = 8'd235;
vramData[13'd385] = 8'd119;
vramData[13'd386] = 8'd176;
vramData[13'd387] = 8'd119;
vramData[13'd388] = 8'd44;
vramData[13'd389] = 8'd247;
vramData[13'd390] = 8'd200;
vramData[13'd391] = 8'd247;
vramData[13'd392] = 8'd16;
vramData[13'd393] = 8'd247;
vramData[13'd394] = 8'd94;
vramData[13'd395] = 8'd55;
vramData[13'd396] = 8'd210;
vramData[13'd397] = 8'd247;
vramData[13'd398] = 8'd16;
vramData[13'd399] = 8'd247;
vramData[13'd400] = 8'd94;
vramData[13'd401] = 8'd135;
vramData[13'd402] = 8'd94;
vramData[13'd403] = 8'd135;
vramData[13'd404] = 8'd223;
vramData[13'd405] = 8'd135;
vramData[13'd406] = 8'd16;
vramData[13'd407] = 8'd120;
vramData[13'd408] = 8'd95;
vramData[13'd409] = 8'd120;
vramData[13'd410] = 8'd95;
vramData[13'd411] = 8'd152;
vramData[13'd412] = 8'd95;
vramData[13'd413] = 8'd152;
vramData[13'd414] = 8'd218;
vramData[13'd415] = 8'd120;
vramData[13'd416] = 8'd223;
vramData[13'd417] = 8'd135;
vramData[13'd418] = 8'd95;
vramData[13'd419] = 8'd120;
vramData[13'd420] = 8'd230;
vramData[13'd421] = 8'd120;
vramData[13'd422] = 8'd6;
vramData[13'd423] = 8'd136;
vramData[13'd424] = 8'd219;
vramData[13'd425] = 8'd129;
vramData[13'd426] = 8'd182;
vramData[13'd427] = 8'd136;
vramData[13'd428] = 8'd183;
vramData[13'd429] = 8'd152;
vramData[13'd430] = 8'd218;
vramData[13'd431] = 8'd120;
vramData[13'd432] = 8'd210;
vramData[13'd433] = 8'd120;
vramData[13'd434] = 8'd30;
vramData[13'd435] = 8'd120;
vramData[13'd436] = 8'd223;
vramData[13'd437] = 8'd120;
vramData[13'd438] = 8'd248;
vramData[13'd439] = 8'd120;
vramData[13'd440] = 8'd165;
vramData[13'd441] = 8'd136;
vramData[13'd442] = 8'd244;
vramData[13'd443] = 8'd136;
vramData[13'd444] = 8'd214;
vramData[13'd445] = 8'd152;
vramData[13'd446] = 8'd30;
vramData[13'd447] = 8'd120;
vramData[13'd448] = 8'd207;
vramData[13'd449] = 8'd120;
vramData[13'd450] = 8'd31;
vramData[13'd451] = 8'd120;
vramData[13'd452] = 8'd30;
vramData[13'd453] = 8'd120;
vramData[13'd454] = 8'd183;
vramData[13'd455] = 8'd120;
vramData[13'd456] = 8'd198;
vramData[13'd457] = 8'd120;
vramData[13'd458] = 8'd135;
vramData[13'd459] = 8'd135;
vramData[13'd460] = 8'd52;
vramData[13'd461] = 8'd87;
vramData[13'd462] = 8'd70;
vramData[13'd463] = 8'd87;
vramData[13'd464] = 8'd39;
vramData[13'd465] = 8'd247;
vramData[13'd466] = 8'd16;
vramData[13'd467] = 8'd247;
vramData[13'd468] = 8'd146;
vramData[13'd469] = 8'd119;
vramData[13'd470] = 8'd255;
vramData[13'd471] = 8'd199;
vramData[13'd472] = 8'd210;
vramData[13'd473] = 8'd55;
vramData[13'd474] = 8'd210;
vramData[13'd475] = 8'd55;
vramData[13'd476] = 8'd164;
vramData[13'd477] = 8'd152;
vramData[13'd478] = 8'd16;
vramData[13'd479] = 8'd135;
vramData[13'd480] = 8'd210;
vramData[13'd481] = 8'd55;
vramData[13'd482] = 8'd202;
vramData[13'd483] = 8'd183;
vramData[13'd484] = 8'd202;
vramData[13'd485] = 8'd183;
vramData[13'd486] = 8'd202;
vramData[13'd487] = 8'd183;
vramData[13'd488] = 8'd202;
vramData[13'd489] = 8'd183;
vramData[13'd490] = 8'd202;
vramData[13'd491] = 8'd183;
vramData[13'd492] = 8'd202;
vramData[13'd493] = 8'd183;
vramData[13'd494] = 8'd202;
vramData[13'd495] = 8'd183;
vramData[13'd496] = 8'd202;
vramData[13'd497] = 8'd183;
vramData[13'd498] = 8'd202;
vramData[13'd499] = 8'd183;
vramData[13'd500] = 8'd31;
vramData[13'd501] = 8'd183;
vramData[13'd502] = 8'd31;
vramData[13'd503] = 8'd183;
vramData[13'd504] = 8'd48;
vramData[13'd505] = 8'd183;
vramData[13'd506] = 8'd37;
vramData[13'd507] = 8'd183;
vramData[13'd508] = 8'd202;
vramData[13'd509] = 8'd183;
vramData[13'd510] = 8'd202;
vramData[13'd511] = 8'd183;
vramData[13'd512] = 8'd202;
vramData[13'd513] = 8'd183;
vramData[13'd514] = 8'd202;
vramData[13'd515] = 8'd183;
vramData[13'd516] = 8'd202;
vramData[13'd517] = 8'd183;
vramData[13'd518] = 8'd202;
vramData[13'd519] = 8'd183;
vramData[13'd520] = 8'd16;
vramData[13'd521] = 8'd183;
vramData[13'd522] = 8'd16;
vramData[13'd523] = 8'd247;
vramData[13'd524] = 8'd16;
vramData[13'd525] = 8'd183;
vramData[13'd526] = 8'd181;
vramData[13'd527] = 8'd135;
vramData[13'd528] = 8'd188;
vramData[13'd529] = 8'd135;
vramData[13'd530] = 8'd252;
vramData[13'd531] = 8'd135;
vramData[13'd532] = 8'd248;
vramData[13'd533] = 8'd55;
vramData[13'd534] = 8'd249;
vramData[13'd535] = 8'd247;
vramData[13'd536] = 8'd40;
vramData[13'd537] = 8'd119;
vramData[13'd538] = 8'd95;
vramData[13'd539] = 8'd55;
vramData[13'd540] = 8'd214;
vramData[13'd541] = 8'd55;
vramData[13'd542] = 8'd183;
vramData[13'd543] = 8'd55;
vramData[13'd544] = 8'd44;
vramData[13'd545] = 8'd87;
vramData[13'd546] = 8'd7;
vramData[13'd547] = 8'd87;
vramData[13'd548] = 8'd97;
vramData[13'd549] = 8'd119;
vramData[13'd550] = 8'd95;
vramData[13'd551] = 8'd55;
vramData[13'd552] = 8'd39;
vramData[13'd553] = 8'd247;
vramData[13'd554] = 8'd32;
vramData[13'd555] = 8'd183;
vramData[13'd556] = 8'd16;
vramData[13'd557] = 8'd247;
vramData[13'd558] = 8'd170;
vramData[13'd559] = 8'd247;
vramData[13'd560] = 8'd249;
vramData[13'd561] = 8'd87;
vramData[13'd562] = 8'd217;
vramData[13'd563] = 8'd247;
vramData[13'd564] = 8'd209;
vramData[13'd565] = 8'd247;
vramData[13'd566] = 8'd106;
vramData[13'd567] = 8'd247;
vramData[13'd568] = 8'd31;
vramData[13'd569] = 8'd247;
vramData[13'd570] = 8'd94;
vramData[13'd571] = 8'd55;
vramData[13'd572] = 8'd17;
vramData[13'd573] = 8'd247;
vramData[13'd574] = 8'd17;
vramData[13'd575] = 8'd247;
vramData[13'd576] = 8'd202;
vramData[13'd577] = 8'd247;
vramData[13'd578] = 8'd7;
vramData[13'd579] = 8'd247;
vramData[13'd580] = 8'd117;
vramData[13'd581] = 8'd247;
vramData[13'd582] = 8'd200;
vramData[13'd583] = 8'd135;
vramData[13'd584] = 8'd220;
vramData[13'd585] = 8'd120;
vramData[13'd586] = 8'd223;
vramData[13'd587] = 8'd135;
vramData[13'd588] = 8'd95;
vramData[13'd589] = 8'd135;
vramData[13'd590] = 8'd210;
vramData[13'd591] = 8'd135;
vramData[13'd592] = 8'd188;
vramData[13'd593] = 8'd120;
vramData[13'd594] = 8'd150;
vramData[13'd595] = 8'd152;
vramData[13'd596] = 8'd16;
vramData[13'd597] = 8'd152;
vramData[13'd598] = 8'd183;
vramData[13'd599] = 8'd136;
vramData[13'd600] = 8'd46;
vramData[13'd601] = 8'd152;
vramData[13'd602] = 8'd214;
vramData[13'd603] = 8'd152;
vramData[13'd604] = 8'd200;
vramData[13'd605] = 8'd120;
vramData[13'd606] = 8'd80;
vramData[13'd607] = 8'd120;
vramData[13'd608] = 8'd55;
vramData[13'd609] = 8'd120;
vramData[13'd610] = 8'd126;
vramData[13'd611] = 8'd120;
vramData[13'd612] = 8'd202;
vramData[13'd613] = 8'd120;
vramData[13'd614] = 8'd31;
vramData[13'd615] = 8'd120;
vramData[13'd616] = 8'd202;
vramData[13'd617] = 8'd135;
vramData[13'd618] = 8'd202;
vramData[13'd619] = 8'd135;
vramData[13'd620] = 8'd16;
vramData[13'd621] = 8'd87;
vramData[13'd622] = 8'd31;
vramData[13'd623] = 8'd247;
vramData[13'd624] = 8'd230;
vramData[13'd625] = 8'd247;
vramData[13'd626] = 8'd156;
vramData[13'd627] = 8'd247;
vramData[13'd628] = 8'd65;
vramData[13'd629] = 8'd119;
vramData[13'd630] = 8'd214;
vramData[13'd631] = 8'd55;
vramData[13'd632] = 8'd210;
vramData[13'd633] = 8'd55;
vramData[13'd634] = 8'd214;
vramData[13'd635] = 8'd135;
vramData[13'd636] = 8'd164;
vramData[13'd637] = 8'd120;
vramData[13'd638] = 8'd16;
vramData[13'd639] = 8'd127;
vramData[13'd640] = 8'd16;
vramData[13'd641] = 8'd8;
vramData[13'd642] = 8'd230;
vramData[13'd643] = 8'd135;
vramData[13'd644] = 8'd31;
vramData[13'd645] = 8'd247;
vramData[13'd646] = 8'd31;
vramData[13'd647] = 8'd247;
vramData[13'd648] = 8'd31;
vramData[13'd649] = 8'd247;
vramData[13'd650] = 8'd30;
vramData[13'd651] = 8'd247;
vramData[13'd652] = 8'd30;
vramData[13'd653] = 8'd247;
vramData[13'd654] = 8'd30;
vramData[13'd655] = 8'd247;
vramData[13'd656] = 8'd30;
vramData[13'd657] = 8'd247;
vramData[13'd658] = 8'd30;
vramData[13'd659] = 8'd247;
vramData[13'd660] = 8'd30;
vramData[13'd661] = 8'd247;
vramData[13'd662] = 8'd210;
vramData[13'd663] = 8'd247;
vramData[13'd664] = 8'd183;
vramData[13'd665] = 8'd247;
vramData[13'd666] = 8'd183;
vramData[13'd667] = 8'd247;
vramData[13'd668] = 8'd252;
vramData[13'd669] = 8'd55;
vramData[13'd670] = 8'd252;
vramData[13'd671] = 8'd55;
vramData[13'd672] = 8'd252;
vramData[13'd673] = 8'd55;
vramData[13'd674] = 8'd252;
vramData[13'd675] = 8'd55;
vramData[13'd676] = 8'd166;
vramData[13'd677] = 8'd55;
vramData[13'd678] = 8'd126;
vramData[13'd679] = 8'd55;
vramData[13'd680] = 8'd39;
vramData[13'd681] = 8'd55;
vramData[13'd682] = 8'd94;
vramData[13'd683] = 8'd247;
vramData[13'd684] = 8'd237;
vramData[13'd685] = 8'd119;
vramData[13'd686] = 8'd210;
vramData[13'd687] = 8'd55;
vramData[13'd688] = 8'd230;
vramData[13'd689] = 8'd135;
vramData[13'd690] = 8'd249;
vramData[13'd691] = 8'd55;
vramData[13'd692] = 8'd213;
vramData[13'd693] = 8'd55;
vramData[13'd694] = 8'd230;
vramData[13'd695] = 8'd135;
vramData[13'd696] = 8'd198;
vramData[13'd697] = 8'd135;
vramData[13'd698] = 8'd198;
vramData[13'd699] = 8'd135;
vramData[13'd700] = 8'd16;
vramData[13'd701] = 8'd135;
vramData[13'd702] = 8'd230;
vramData[13'd703] = 8'd135;
vramData[13'd704] = 8'd230;
vramData[13'd705] = 8'd135;
vramData[13'd706] = 8'd19;
vramData[13'd707] = 8'd135;
vramData[13'd708] = 8'd17;
vramData[13'd709] = 8'd55;
vramData[13'd710] = 8'd96;
vramData[13'd711] = 8'd55;
vramData[13'd712] = 8'd0;
vramData[13'd713] = 8'd71;
vramData[13'd714] = 8'd44;
vramData[13'd715] = 8'd135;
vramData[13'd716] = 8'd96;
vramData[13'd717] = 8'd247;
vramData[13'd718] = 8'd251;
vramData[13'd719] = 8'd247;
vramData[13'd720] = 8'd212;
vramData[13'd721] = 8'd247;
vramData[13'd722] = 8'd44;
vramData[13'd723] = 8'd247;
vramData[13'd724] = 8'd249;
vramData[13'd725] = 8'd55;
vramData[13'd726] = 8'd7;
vramData[13'd727] = 8'd55;
vramData[13'd728] = 8'd250;
vramData[13'd729] = 8'd247;
vramData[13'd730] = 8'd166;
vramData[13'd731] = 8'd55;
vramData[13'd732] = 8'd135;
vramData[13'd733] = 8'd247;
vramData[13'd734] = 8'd44;
vramData[13'd735] = 8'd103;
vramData[13'd736] = 8'd192;
vramData[13'd737] = 8'd135;
vramData[13'd738] = 8'd17;
vramData[13'd739] = 8'd135;
vramData[13'd740] = 8'd214;
vramData[13'd741] = 8'd135;
vramData[13'd742] = 8'd16;
vramData[13'd743] = 8'd135;
vramData[13'd744] = 8'd183;
vramData[13'd745] = 8'd135;
vramData[13'd746] = 8'd214;
vramData[13'd747] = 8'd135;
vramData[13'd748] = 8'd148;
vramData[13'd749] = 8'd120;
vramData[13'd750] = 8'd16;
vramData[13'd751] = 8'd120;
vramData[13'd752] = 8'd135;
vramData[13'd753] = 8'd120;
vramData[13'd754] = 8'd230;
vramData[13'd755] = 8'd120;
vramData[13'd756] = 8'd76;
vramData[13'd757] = 8'd120;
vramData[13'd758] = 8'd95;
vramData[13'd759] = 8'd120;
vramData[13'd760] = 8'd31;
vramData[13'd761] = 8'd152;
vramData[13'd762] = 8'd102;
vramData[13'd763] = 8'd120;
vramData[13'd764] = 8'd9;
vramData[13'd765] = 8'd120;
vramData[13'd766] = 8'd202;
vramData[13'd767] = 8'd120;
vramData[13'd768] = 8'd31;
vramData[13'd769] = 8'd120;
vramData[13'd770] = 8'd202;
vramData[13'd771] = 8'd120;
vramData[13'd772] = 8'd164;
vramData[13'd773] = 8'd135;
vramData[13'd774] = 8'd230;
vramData[13'd775] = 8'd135;
vramData[13'd776] = 8'd126;
vramData[13'd777] = 8'd135;
vramData[13'd778] = 8'd167;
vramData[13'd779] = 8'd135;
vramData[13'd780] = 8'd46;
vramData[13'd781] = 8'd135;
vramData[13'd782] = 8'd214;
vramData[13'd783] = 8'd247;
vramData[13'd784] = 8'd253;
vramData[13'd785] = 8'd247;
vramData[13'd786] = 8'd96;
vramData[13'd787] = 8'd247;
vramData[13'd788] = 8'd214;
vramData[13'd789] = 8'd55;
vramData[13'd790] = 8'd210;
vramData[13'd791] = 8'd55;
vramData[13'd792] = 8'd210;
vramData[13'd793] = 8'd55;
vramData[13'd794] = 8'd16;
vramData[13'd795] = 8'd120;
vramData[13'd796] = 8'd221;
vramData[13'd797] = 8'd135;
vramData[13'd798] = 8'd85;
vramData[13'd799] = 8'd127;
vramData[13'd800] = 8'd202;
vramData[13'd801] = 8'd8;
vramData[13'd802] = 8'd16;
vramData[13'd803] = 8'd8;
vramData[13'd804] = 8'd16;
vramData[13'd805] = 8'd135;
vramData[13'd806] = 8'd16;
vramData[13'd807] = 8'd103;
vramData[13'd808] = 8'd16;
vramData[13'd809] = 8'd103;
vramData[13'd810] = 8'd30;
vramData[13'd811] = 8'd103;
vramData[13'd812] = 8'd16;
vramData[13'd813] = 8'd103;
vramData[13'd814] = 8'd164;
vramData[13'd815] = 8'd103;
vramData[13'd816] = 8'd209;
vramData[13'd817] = 8'd231;
vramData[13'd818] = 8'd210;
vramData[13'd819] = 8'd247;
vramData[13'd820] = 8'd210;
vramData[13'd821] = 8'd247;
vramData[13'd822] = 8'd210;
vramData[13'd823] = 8'd247;
vramData[13'd824] = 8'd210;
vramData[13'd825] = 8'd247;
vramData[13'd826] = 8'd30;
vramData[13'd827] = 8'd247;
vramData[13'd828] = 8'd95;
vramData[13'd829] = 8'd247;
vramData[13'd830] = 8'd250;
vramData[13'd831] = 8'd247;
vramData[13'd832] = 8'd94;
vramData[13'd833] = 8'd247;
vramData[13'd834] = 8'd94;
vramData[13'd835] = 8'd247;
vramData[13'd836] = 8'd189;
vramData[13'd837] = 8'd119;
vramData[13'd838] = 8'd95;
vramData[13'd839] = 8'd55;
vramData[13'd840] = 8'd210;
vramData[13'd841] = 8'd55;
vramData[13'd842] = 8'd214;
vramData[13'd843] = 8'd135;
vramData[13'd844] = 8'd210;
vramData[13'd845] = 8'd135;
vramData[13'd846] = 8'd198;
vramData[13'd847] = 8'd135;
vramData[13'd848] = 8'd16;
vramData[13'd849] = 8'd135;
vramData[13'd850] = 8'd16;
vramData[13'd851] = 8'd135;
vramData[13'd852] = 8'd80;
vramData[13'd853] = 8'd120;
vramData[13'd854] = 8'd202;
vramData[13'd855] = 8'd120;
vramData[13'd856] = 8'd16;
vramData[13'd857] = 8'd135;
vramData[13'd858] = 8'd159;
vramData[13'd859] = 8'd135;
vramData[13'd860] = 8'd16;
vramData[13'd861] = 8'd120;
vramData[13'd862] = 8'd135;
vramData[13'd863] = 8'd135;
vramData[13'd864] = 8'd37;
vramData[13'd865] = 8'd135;
vramData[13'd866] = 8'd17;
vramData[13'd867] = 8'd135;
vramData[13'd868] = 8'd53;
vramData[13'd869] = 8'd119;
vramData[13'd870] = 8'd179;
vramData[13'd871] = 8'd87;
vramData[13'd872] = 8'd95;
vramData[13'd873] = 8'd87;
vramData[13'd874] = 8'd96;
vramData[13'd875] = 8'd135;
vramData[13'd876] = 8'd214;
vramData[13'd877] = 8'd247;
vramData[13'd878] = 8'd183;
vramData[13'd879] = 8'd103;
vramData[13'd880] = 8'd126;
vramData[13'd881] = 8'd247;
vramData[13'd882] = 8'd94;
vramData[13'd883] = 8'd247;
vramData[13'd884] = 8'd226;
vramData[13'd885] = 8'd247;
vramData[13'd886] = 8'd39;
vramData[13'd887] = 8'd247;
vramData[13'd888] = 8'd152;
vramData[13'd889] = 8'd119;
vramData[13'd890] = 8'd39;
vramData[13'd891] = 8'd247;
vramData[13'd892] = 8'd44;
vramData[13'd893] = 8'd135;
vramData[13'd894] = 8'd189;
vramData[13'd895] = 8'd103;
vramData[13'd896] = 8'd95;
vramData[13'd897] = 8'd135;
vramData[13'd898] = 8'd90;
vramData[13'd899] = 8'd135;
vramData[13'd900] = 8'd202;
vramData[13'd901] = 8'd135;
vramData[13'd902] = 8'd17;
vramData[13'd903] = 8'd120;
vramData[13'd904] = 8'd85;
vramData[13'd905] = 8'd135;
vramData[13'd906] = 8'd16;
vramData[13'd907] = 8'd120;
vramData[13'd908] = 8'd210;
vramData[13'd909] = 8'd120;
vramData[13'd910] = 8'd188;
vramData[13'd911] = 8'd120;
vramData[13'd912] = 8'd202;
vramData[13'd913] = 8'd120;
vramData[13'd914] = 8'd253;
vramData[13'd915] = 8'd120;
vramData[13'd916] = 8'd198;
vramData[13'd917] = 8'd120;
vramData[13'd918] = 8'd198;
vramData[13'd919] = 8'd120;
vramData[13'd920] = 8'd230;
vramData[13'd921] = 8'd120;
vramData[13'd922] = 8'd16;
vramData[13'd923] = 8'd120;
vramData[13'd924] = 8'd9;
vramData[13'd925] = 8'd120;
vramData[13'd926] = 8'd31;
vramData[13'd927] = 8'd120;
vramData[13'd928] = 8'd37;
vramData[13'd929] = 8'd120;
vramData[13'd930] = 8'd85;
vramData[13'd931] = 8'd120;
vramData[13'd932] = 8'd37;
vramData[13'd933] = 8'd120;
vramData[13'd934] = 8'd210;
vramData[13'd935] = 8'd135;
vramData[13'd936] = 8'd183;
vramData[13'd937] = 8'd135;
vramData[13'd938] = 8'd17;
vramData[13'd939] = 8'd135;
vramData[13'd940] = 8'd29;
vramData[13'd941] = 8'd247;
vramData[13'd942] = 8'd229;
vramData[13'd943] = 8'd247;
vramData[13'd944] = 8'd46;
vramData[13'd945] = 8'd247;
vramData[13'd946] = 8'd210;
vramData[13'd947] = 8'd55;
vramData[13'd948] = 8'd210;
vramData[13'd949] = 8'd135;
vramData[13'd950] = 8'd210;
vramData[13'd951] = 8'd135;
vramData[13'd952] = 8'd210;
vramData[13'd953] = 8'd135;
vramData[13'd954] = 8'd70;
vramData[13'd955] = 8'd120;
vramData[13'd956] = 8'd16;
vramData[13'd957] = 8'd135;
vramData[13'd958] = 8'd80;
vramData[13'd959] = 8'd123;
vramData[13'd960] = 8'd210;
vramData[13'd961] = 8'd8;
vramData[13'd962] = 8'd65;
vramData[13'd963] = 8'd136;
vramData[13'd964] = 8'd135;
vramData[13'd965] = 8'd135;
vramData[13'd966] = 8'd210;
vramData[13'd967] = 8'd103;
vramData[13'd968] = 8'd210;
vramData[13'd969] = 8'd103;
vramData[13'd970] = 8'd210;
vramData[13'd971] = 8'd103;
vramData[13'd972] = 8'd210;
vramData[13'd973] = 8'd103;
vramData[13'd974] = 8'd183;
vramData[13'd975] = 8'd103;
vramData[13'd976] = 8'd202;
vramData[13'd977] = 8'd231;
vramData[13'd978] = 8'd30;
vramData[13'd979] = 8'd247;
vramData[13'd980] = 8'd30;
vramData[13'd981] = 8'd247;
vramData[13'd982] = 8'd30;
vramData[13'd983] = 8'd247;
vramData[13'd984] = 8'd16;
vramData[13'd985] = 8'd247;
vramData[13'd986] = 8'd16;
vramData[13'd987] = 8'd247;
vramData[13'd988] = 8'd45;
vramData[13'd989] = 8'd247;
vramData[13'd990] = 8'd95;
vramData[13'd991] = 8'd135;
vramData[13'd992] = 8'd183;
vramData[13'd993] = 8'd135;
vramData[13'd994] = 8'd209;
vramData[13'd995] = 8'd135;
vramData[13'd996] = 8'd210;
vramData[13'd997] = 8'd135;
vramData[13'd998] = 8'd202;
vramData[13'd999] = 8'd120;
vramData[13'd1000] = 8'd80;
vramData[13'd1001] = 8'd120;
vramData[13'd1002] = 8'd202;
vramData[13'd1003] = 8'd152;
vramData[13'd1004] = 8'd198;
vramData[13'd1005] = 8'd152;
vramData[13'd1006] = 8'd200;
vramData[13'd1007] = 8'd120;
vramData[13'd1008] = 8'd181;
vramData[13'd1009] = 8'd120;
vramData[13'd1010] = 8'd85;
vramData[13'd1011] = 8'd120;
vramData[13'd1012] = 8'd181;
vramData[13'd1013] = 8'd135;
vramData[13'd1014] = 8'd135;
vramData[13'd1015] = 8'd120;
vramData[13'd1016] = 8'd208;
vramData[13'd1017] = 8'd120;
vramData[13'd1018] = 8'd188;
vramData[13'd1019] = 8'd120;
vramData[13'd1020] = 8'd30;
vramData[13'd1021] = 8'd120;
vramData[13'd1022] = 8'd164;
vramData[13'd1023] = 8'd120;
vramData[13'd1024] = 8'd148;
vramData[13'd1025] = 8'd135;
vramData[13'd1026] = 8'd17;
vramData[13'd1027] = 8'd135;
vramData[13'd1028] = 8'd209;
vramData[13'd1029] = 8'd55;
vramData[13'd1030] = 8'd198;
vramData[13'd1031] = 8'd135;
vramData[13'd1032] = 8'd16;
vramData[13'd1033] = 8'd135;
vramData[13'd1034] = 8'd95;
vramData[13'd1035] = 8'd135;
vramData[13'd1036] = 8'd12;
vramData[13'd1037] = 8'd119;
vramData[13'd1038] = 8'd180;
vramData[13'd1039] = 8'd87;
vramData[13'd1040] = 8'd183;
vramData[13'd1041] = 8'd103;
vramData[13'd1042] = 8'd7;
vramData[13'd1043] = 8'd135;
vramData[13'd1044] = 8'd213;
vramData[13'd1045] = 8'd55;
vramData[13'd1046] = 8'd210;
vramData[13'd1047] = 8'd135;
vramData[13'd1048] = 8'd85;
vramData[13'd1049] = 8'd120;
vramData[13'd1050] = 8'd248;
vramData[13'd1051] = 8'd120;
vramData[13'd1052] = 8'd198;
vramData[13'd1053] = 8'd120;
vramData[13'd1054] = 8'd210;
vramData[13'd1055] = 8'd135;
vramData[13'd1056] = 8'd109;
vramData[13'd1057] = 8'd135;
vramData[13'd1058] = 8'd16;
vramData[13'd1059] = 8'd135;
vramData[13'd1060] = 8'd210;
vramData[13'd1061] = 8'd135;
vramData[13'd1062] = 8'd181;
vramData[13'd1063] = 8'd135;
vramData[13'd1064] = 8'd210;
vramData[13'd1065] = 8'd135;
vramData[13'd1066] = 8'd85;
vramData[13'd1067] = 8'd135;
vramData[13'd1068] = 8'd90;
vramData[13'd1069] = 8'd120;
vramData[13'd1070] = 8'd210;
vramData[13'd1071] = 8'd120;
vramData[13'd1072] = 8'd16;
vramData[13'd1073] = 8'd120;
vramData[13'd1074] = 8'd31;
vramData[13'd1075] = 8'd120;
vramData[13'd1076] = 8'd30;
vramData[13'd1077] = 8'd120;
vramData[13'd1078] = 8'd164;
vramData[13'd1079] = 8'd120;
vramData[13'd1080] = 8'd16;
vramData[13'd1081] = 8'd120;
vramData[13'd1082] = 8'd213;
vramData[13'd1083] = 8'd120;
vramData[13'd1084] = 8'd210;
vramData[13'd1085] = 8'd120;
vramData[13'd1086] = 8'd16;
vramData[13'd1087] = 8'd120;
vramData[13'd1088] = 8'd202;
vramData[13'd1089] = 8'd135;
vramData[13'd1090] = 8'd202;
vramData[13'd1091] = 8'd135;
vramData[13'd1092] = 8'd248;
vramData[13'd1093] = 8'd135;
vramData[13'd1094] = 8'd126;
vramData[13'd1095] = 8'd135;
vramData[13'd1096] = 8'd248;
vramData[13'd1097] = 8'd135;
vramData[13'd1098] = 8'd55;
vramData[13'd1099] = 8'd135;
vramData[13'd1100] = 8'd37;
vramData[13'd1101] = 8'd55;
vramData[13'd1102] = 8'd31;
vramData[13'd1103] = 8'd135;
vramData[13'd1104] = 8'd34;
vramData[13'd1105] = 8'd247;
vramData[13'd1106] = 8'd200;
vramData[13'd1107] = 8'd55;
vramData[13'd1108] = 8'd202;
vramData[13'd1109] = 8'd55;
vramData[13'd1110] = 8'd83;
vramData[13'd1111] = 8'd135;
vramData[13'd1112] = 8'd80;
vramData[13'd1113] = 8'd120;
vramData[13'd1114] = 8'd210;
vramData[13'd1115] = 8'd120;
vramData[13'd1116] = 8'd210;
vramData[13'd1117] = 8'd55;
vramData[13'd1118] = 8'd202;
vramData[13'd1119] = 8'd179;
vramData[13'd1120] = 8'd16;
vramData[13'd1121] = 8'd24;
vramData[13'd1122] = 8'd214;
vramData[13'd1123] = 8'd120;
vramData[13'd1124] = 8'd220;
vramData[13'd1125] = 8'd120;
vramData[13'd1126] = 8'd220;
vramData[13'd1127] = 8'd120;
vramData[13'd1128] = 8'd223;
vramData[13'd1129] = 8'd135;
vramData[13'd1130] = 8'd223;
vramData[13'd1131] = 8'd135;
vramData[13'd1132] = 8'd223;
vramData[13'd1133] = 8'd135;
vramData[13'd1134] = 8'd220;
vramData[13'd1135] = 8'd120;
vramData[13'd1136] = 8'd223;
vramData[13'd1137] = 8'd135;
vramData[13'd1138] = 8'd31;
vramData[13'd1139] = 8'd135;
vramData[13'd1140] = 8'd31;
vramData[13'd1141] = 8'd135;
vramData[13'd1142] = 8'd31;
vramData[13'd1143] = 8'd135;
vramData[13'd1144] = 8'd31;
vramData[13'd1145] = 8'd135;
vramData[13'd1146] = 8'd30;
vramData[13'd1147] = 8'd135;
vramData[13'd1148] = 8'd210;
vramData[13'd1149] = 8'd135;
vramData[13'd1150] = 8'd202;
vramData[13'd1151] = 8'd120;
vramData[13'd1152] = 8'd248;
vramData[13'd1153] = 8'd120;
vramData[13'd1154] = 8'd94;
vramData[13'd1155] = 8'd120;
vramData[13'd1156] = 8'd211;
vramData[13'd1157] = 8'd120;
vramData[13'd1158] = 8'd16;
vramData[13'd1159] = 8'd120;
vramData[13'd1160] = 8'd94;
vramData[13'd1161] = 8'd152;
vramData[13'd1162] = 8'd94;
vramData[13'd1163] = 8'd8;
vramData[13'd1164] = 8'd212;
vramData[13'd1165] = 8'd152;
vramData[13'd1166] = 8'd181;
vramData[13'd1167] = 8'd152;
vramData[13'd1168] = 8'd202;
vramData[13'd1169] = 8'd152;
vramData[13'd1170] = 8'd166;
vramData[13'd1171] = 8'd120;
vramData[13'd1172] = 8'd210;
vramData[13'd1173] = 8'd120;
vramData[13'd1174] = 8'd85;
vramData[13'd1175] = 8'd120;
vramData[13'd1176] = 8'd148;
vramData[13'd1177] = 8'd120;
vramData[13'd1178] = 8'd230;
vramData[13'd1179] = 8'd120;
vramData[13'd1180] = 8'd164;
vramData[13'd1181] = 8'd152;
vramData[13'd1182] = 8'd194;
vramData[13'd1183] = 8'd120;
vramData[13'd1184] = 8'd80;
vramData[13'd1185] = 8'd135;
vramData[13'd1186] = 8'd181;
vramData[13'd1187] = 8'd135;
vramData[13'd1188] = 8'd16;
vramData[13'd1189] = 8'd135;
vramData[13'd1190] = 8'd31;
vramData[13'd1191] = 8'd135;
vramData[13'd1192] = 8'd164;
vramData[13'd1193] = 8'd135;
vramData[13'd1194] = 8'd218;
vramData[13'd1195] = 8'd135;
vramData[13'd1196] = 8'd184;
vramData[13'd1197] = 8'd135;
vramData[13'd1198] = 8'd95;
vramData[13'd1199] = 8'd87;
vramData[13'd1200] = 8'd95;
vramData[13'd1201] = 8'd135;
vramData[13'd1202] = 8'd202;
vramData[13'd1203] = 8'd120;
vramData[13'd1204] = 8'd80;
vramData[13'd1205] = 8'd120;
vramData[13'd1206] = 8'd252;
vramData[13'd1207] = 8'd120;
vramData[13'd1208] = 8'd202;
vramData[13'd1209] = 8'd120;
vramData[13'd1210] = 8'd85;
vramData[13'd1211] = 8'd120;
vramData[13'd1212] = 8'd150;
vramData[13'd1213] = 8'd120;
vramData[13'd1214] = 8'd172;
vramData[13'd1215] = 8'd135;
vramData[13'd1216] = 8'd164;
vramData[13'd1217] = 8'd135;
vramData[13'd1218] = 8'd202;
vramData[13'd1219] = 8'd120;
vramData[13'd1220] = 8'd181;
vramData[13'd1221] = 8'd120;
vramData[13'd1222] = 8'd210;
vramData[13'd1223] = 8'd120;
vramData[13'd1224] = 8'd85;
vramData[13'd1225] = 8'd120;
vramData[13'd1226] = 8'd230;
vramData[13'd1227] = 8'd135;
vramData[13'd1228] = 8'd171;
vramData[13'd1229] = 8'd135;
vramData[13'd1230] = 8'd198;
vramData[13'd1231] = 8'd135;
vramData[13'd1232] = 8'd197;
vramData[13'd1233] = 8'd135;
vramData[13'd1234] = 8'd230;
vramData[13'd1235] = 8'd120;
vramData[13'd1236] = 8'd210;
vramData[13'd1237] = 8'd120;
vramData[13'd1238] = 8'd31;
vramData[13'd1239] = 8'd120;
vramData[13'd1240] = 8'd135;
vramData[13'd1241] = 8'd120;
vramData[13'd1242] = 8'd31;
vramData[13'd1243] = 8'd120;
vramData[13'd1244] = 8'd31;
vramData[13'd1245] = 8'd120;
vramData[13'd1246] = 8'd16;
vramData[13'd1247] = 8'd135;
vramData[13'd1248] = 8'd214;
vramData[13'd1249] = 8'd135;
vramData[13'd1250] = 8'd30;
vramData[13'd1251] = 8'd87;
vramData[13'd1252] = 8'd16;
vramData[13'd1253] = 8'd87;
vramData[13'd1254] = 8'd28;
vramData[13'd1255] = 8'd87;
vramData[13'd1256] = 8'd214;
vramData[13'd1257] = 8'd55;
vramData[13'd1258] = 8'd210;
vramData[13'd1259] = 8'd55;
vramData[13'd1260] = 8'd16;
vramData[13'd1261] = 8'd55;
vramData[13'd1262] = 8'd114;
vramData[13'd1263] = 8'd119;
vramData[13'd1264] = 8'd32;
vramData[13'd1265] = 8'd167;
vramData[13'd1266] = 8'd207;
vramData[13'd1267] = 8'd55;
vramData[13'd1268] = 8'd31;
vramData[13'd1269] = 8'd55;
vramData[13'd1270] = 8'd214;
vramData[13'd1271] = 8'd135;
vramData[13'd1272] = 8'd16;
vramData[13'd1273] = 8'd135;
vramData[13'd1274] = 8'd214;
vramData[13'd1275] = 8'd135;
vramData[13'd1276] = 8'd95;
vramData[13'd1277] = 8'd135;
vramData[13'd1278] = 8'd95;
vramData[13'd1279] = 8'd135;
vramData[13'd1280] = 8'd210;
vramData[13'd1281] = 8'd24;
vramData[13'd1282] = 8'd16;
vramData[13'd1283] = 8'd8;
vramData[13'd1284] = 8'd230;
vramData[13'd1285] = 8'd135;
vramData[13'd1286] = 8'd252;
vramData[13'd1287] = 8'd247;
vramData[13'd1288] = 8'd200;
vramData[13'd1289] = 8'd247;
vramData[13'd1290] = 8'd202;
vramData[13'd1291] = 8'd247;
vramData[13'd1292] = 8'd202;
vramData[13'd1293] = 8'd247;
vramData[13'd1294] = 8'd202;
vramData[13'd1295] = 8'd247;
vramData[13'd1296] = 8'd202;
vramData[13'd1297] = 8'd247;
vramData[13'd1298] = 8'd202;
vramData[13'd1299] = 8'd247;
vramData[13'd1300] = 8'd202;
vramData[13'd1301] = 8'd247;
vramData[13'd1302] = 8'd31;
vramData[13'd1303] = 8'd247;
vramData[13'd1304] = 8'd255;
vramData[13'd1305] = 8'd231;
vramData[13'd1306] = 8'd213;
vramData[13'd1307] = 8'd87;
vramData[13'd1308] = 8'd16;
vramData[13'd1309] = 8'd120;
vramData[13'd1310] = 8'd16;
vramData[13'd1311] = 8'd152;
vramData[13'd1312] = 8'd94;
vramData[13'd1313] = 8'd8;
vramData[13'd1314] = 8'd73;
vramData[13'd1315] = 8'd8;
vramData[13'd1316] = 8'd95;
vramData[13'd1317] = 8'd120;
vramData[13'd1318] = 8'd46;
vramData[13'd1319] = 8'd8;
vramData[13'd1320] = 8'd171;
vramData[13'd1321] = 8'd168;
vramData[13'd1322] = 8'd135;
vramData[13'd1323] = 8'd120;
vramData[13'd1324] = 8'd17;
vramData[13'd1325] = 8'd120;
vramData[13'd1326] = 8'd198;
vramData[13'd1327] = 8'd152;
vramData[13'd1328] = 8'd85;
vramData[13'd1329] = 8'd152;
vramData[13'd1330] = 8'd214;
vramData[13'd1331] = 8'd152;
vramData[13'd1332] = 8'd209;
vramData[13'd1333] = 8'd120;
vramData[13'd1334] = 8'd230;
vramData[13'd1335] = 8'd135;
vramData[13'd1336] = 8'd181;
vramData[13'd1337] = 8'd120;
vramData[13'd1338] = 8'd16;
vramData[13'd1339] = 8'd135;
vramData[13'd1340] = 8'd16;
vramData[13'd1341] = 8'd120;
vramData[13'd1342] = 8'd181;
vramData[13'd1343] = 8'd120;
vramData[13'd1344] = 8'd150;
vramData[13'd1345] = 8'd135;
vramData[13'd1346] = 8'd202;
vramData[13'd1347] = 8'd120;
vramData[13'd1348] = 8'd209;
vramData[13'd1349] = 8'd135;
vramData[13'd1350] = 8'd75;
vramData[13'd1351] = 8'd135;
vramData[13'd1352] = 8'd30;
vramData[13'd1353] = 8'd135;
vramData[13'd1354] = 8'd210;
vramData[13'd1355] = 8'd135;
vramData[13'd1356] = 8'd198;
vramData[13'd1357] = 8'd135;
vramData[13'd1358] = 8'd210;
vramData[13'd1359] = 8'd135;
vramData[13'd1360] = 8'd80;
vramData[13'd1361] = 8'd120;
vramData[13'd1362] = 8'd226;
vramData[13'd1363] = 8'd120;
vramData[13'd1364] = 8'd74;
vramData[13'd1365] = 8'd8;
vramData[13'd1366] = 8'd76;
vramData[13'd1367] = 8'd8;
vramData[13'd1368] = 8'd16;
vramData[13'd1369] = 8'd120;
vramData[13'd1370] = 8'd31;
vramData[13'd1371] = 8'd120;
vramData[13'd1372] = 8'd30;
vramData[13'd1373] = 8'd120;
vramData[13'd1374] = 8'd80;
vramData[13'd1375] = 8'd135;
vramData[13'd1376] = 8'd150;
vramData[13'd1377] = 8'd120;
vramData[13'd1378] = 8'd31;
vramData[13'd1379] = 8'd120;
vramData[13'd1380] = 8'd150;
vramData[13'd1381] = 8'd120;
vramData[13'd1382] = 8'd16;
vramData[13'd1383] = 8'd120;
vramData[13'd1384] = 8'd209;
vramData[13'd1385] = 8'd120;
vramData[13'd1386] = 8'd198;
vramData[13'd1387] = 8'd120;
vramData[13'd1388] = 8'd198;
vramData[13'd1389] = 8'd120;
vramData[13'd1390] = 8'd16;
vramData[13'd1391] = 8'd120;
vramData[13'd1392] = 8'd181;
vramData[13'd1393] = 8'd120;
vramData[13'd1394] = 8'd210;
vramData[13'd1395] = 8'd120;
vramData[13'd1396] = 8'd80;
vramData[13'd1397] = 8'd135;
vramData[13'd1398] = 8'd202;
vramData[13'd1399] = 8'd120;
vramData[13'd1400] = 8'd171;
vramData[13'd1401] = 8'd120;
vramData[13'd1402] = 8'd162;
vramData[13'd1403] = 8'd120;
vramData[13'd1404] = 8'd80;
vramData[13'd1405] = 8'd120;
vramData[13'd1406] = 8'd51;
vramData[13'd1407] = 8'd120;
vramData[13'd1408] = 8'd202;
vramData[13'd1409] = 8'd120;
vramData[13'd1410] = 8'd16;
vramData[13'd1411] = 8'd135;
vramData[13'd1412] = 8'd31;
vramData[13'd1413] = 8'd135;
vramData[13'd1414] = 8'd31;
vramData[13'd1415] = 8'd135;
vramData[13'd1416] = 8'd145;
vramData[13'd1417] = 8'd120;
vramData[13'd1418] = 8'd16;
vramData[13'd1419] = 8'd135;
vramData[13'd1420] = 8'd230;
vramData[13'd1421] = 8'd55;
vramData[13'd1422] = 8'd95;
vramData[13'd1423] = 8'd55;
vramData[13'd1424] = 8'd95;
vramData[13'd1425] = 8'd55;
vramData[13'd1426] = 8'd147;
vramData[13'd1427] = 8'd119;
vramData[13'd1428] = 8'd214;
vramData[13'd1429] = 8'd55;
vramData[13'd1430] = 8'd188;
vramData[13'd1431] = 8'd135;
vramData[13'd1432] = 8'd85;
vramData[13'd1433] = 8'd55;
vramData[13'd1434] = 8'd210;
vramData[13'd1435] = 8'd56;
vramData[13'd1436] = 8'd210;
vramData[13'd1437] = 8'd56;
vramData[13'd1438] = 8'd210;
vramData[13'd1439] = 8'd56;
vramData[13'd1440] = 8'd202;
vramData[13'd1441] = 8'd131;
vramData[13'd1442] = 8'd198;
vramData[13'd1443] = 8'd120;
vramData[13'd1444] = 8'd214;
vramData[13'd1445] = 8'd247;
vramData[13'd1446] = 8'd210;
vramData[13'd1447] = 8'd247;
vramData[13'd1448] = 8'd210;
vramData[13'd1449] = 8'd247;
vramData[13'd1450] = 8'd210;
vramData[13'd1451] = 8'd247;
vramData[13'd1452] = 8'd210;
vramData[13'd1453] = 8'd247;
vramData[13'd1454] = 8'd183;
vramData[13'd1455] = 8'd247;
vramData[13'd1456] = 8'd183;
vramData[13'd1457] = 8'd247;
vramData[13'd1458] = 8'd95;
vramData[13'd1459] = 8'd247;
vramData[13'd1460] = 8'd248;
vramData[13'd1461] = 8'd135;
vramData[13'd1462] = 8'd252;
vramData[13'd1463] = 8'd135;
vramData[13'd1464] = 8'd31;
vramData[13'd1465] = 8'd135;
vramData[13'd1466] = 8'd31;
vramData[13'd1467] = 8'd135;
vramData[13'd1468] = 8'd16;
vramData[13'd1469] = 8'd120;
vramData[13'd1470] = 8'd226;
vramData[13'd1471] = 8'd200;
vramData[13'd1472] = 8'd214;
vramData[13'd1473] = 8'd120;
vramData[13'd1474] = 8'd202;
vramData[13'd1475] = 8'd55;
vramData[13'd1476] = 8'd164;
vramData[13'd1477] = 8'd115;
vramData[13'd1478] = 8'd16;
vramData[13'd1479] = 8'd56;
vramData[13'd1480] = 8'd31;
vramData[13'd1481] = 8'd56;
vramData[13'd1482] = 8'd135;
vramData[13'd1483] = 8'd120;
vramData[13'd1484] = 8'd30;
vramData[13'd1485] = 8'd120;
vramData[13'd1486] = 8'd209;
vramData[13'd1487] = 8'd120;
vramData[13'd1488] = 8'd210;
vramData[13'd1489] = 8'd152;
vramData[13'd1490] = 8'd210;
vramData[13'd1491] = 8'd120;
vramData[13'd1492] = 8'd202;
vramData[13'd1493] = 8'd135;
vramData[13'd1494] = 8'd16;
vramData[13'd1495] = 8'd135;
vramData[13'd1496] = 8'd164;
vramData[13'd1497] = 8'd135;
vramData[13'd1498] = 8'd16;
vramData[13'd1499] = 8'd135;
vramData[13'd1500] = 8'd164;
vramData[13'd1501] = 8'd135;
vramData[13'd1502] = 8'd214;
vramData[13'd1503] = 8'd135;
vramData[13'd1504] = 8'd212;
vramData[13'd1505] = 8'd135;
vramData[13'd1506] = 8'd17;
vramData[13'd1507] = 8'd120;
vramData[13'd1508] = 8'd188;
vramData[13'd1509] = 8'd120;
vramData[13'd1510] = 8'd200;
vramData[13'd1511] = 8'd120;
vramData[13'd1512] = 8'd31;
vramData[13'd1513] = 8'd120;
vramData[13'd1514] = 8'd30;
vramData[13'd1515] = 8'd120;
vramData[13'd1516] = 8'd17;
vramData[13'd1517] = 8'd135;
vramData[13'd1518] = 8'd31;
vramData[13'd1519] = 8'd120;
vramData[13'd1520] = 8'd213;
vramData[13'd1521] = 8'd8;
vramData[13'd1522] = 8'd16;
vramData[13'd1523] = 8'd8;
vramData[13'd1524] = 8'd110;
vramData[13'd1525] = 8'd8;
vramData[13'd1526] = 8'd44;
vramData[13'd1527] = 8'd120;
vramData[13'd1528] = 8'd214;
vramData[13'd1529] = 8'd120;
vramData[13'd1530] = 8'd85;
vramData[13'd1531] = 8'd120;
vramData[13'd1532] = 8'd166;
vramData[13'd1533] = 8'd120;
vramData[13'd1534] = 8'd80;
vramData[13'd1535] = 8'd120;
vramData[13'd1536] = 8'd31;
vramData[13'd1537] = 8'd120;
vramData[13'd1538] = 8'd202;
vramData[13'd1539] = 8'd120;
vramData[13'd1540] = 8'd230;
vramData[13'd1541] = 8'd120;
vramData[13'd1542] = 8'd17;
vramData[13'd1543] = 8'd120;
vramData[13'd1544] = 8'd37;
vramData[13'd1545] = 8'd135;
vramData[13'd1546] = 8'd16;
vramData[13'd1547] = 8'd120;
vramData[13'd1548] = 8'd181;
vramData[13'd1549] = 8'd120;
vramData[13'd1550] = 8'd135;
vramData[13'd1551] = 8'd120;
vramData[13'd1552] = 8'd202;
vramData[13'd1553] = 8'd120;
vramData[13'd1554] = 8'd16;
vramData[13'd1555] = 8'd135;
vramData[13'd1556] = 8'd30;
vramData[13'd1557] = 8'd135;
vramData[13'd1558] = 8'd210;
vramData[13'd1559] = 8'd120;
vramData[13'd1560] = 8'd135;
vramData[13'd1561] = 8'd120;
vramData[13'd1562] = 8'd135;
vramData[13'd1563] = 8'd120;
vramData[13'd1564] = 8'd16;
vramData[13'd1565] = 8'd120;
vramData[13'd1566] = 8'd16;
vramData[13'd1567] = 8'd120;
vramData[13'd1568] = 8'd135;
vramData[13'd1569] = 8'd120;
vramData[13'd1570] = 8'd31;
vramData[13'd1571] = 8'd120;
vramData[13'd1572] = 8'd202;
vramData[13'd1573] = 8'd120;
vramData[13'd1574] = 8'd16;
vramData[13'd1575] = 8'd135;
vramData[13'd1576] = 8'd16;
vramData[13'd1577] = 8'd120;
vramData[13'd1578] = 8'd83;
vramData[13'd1579] = 8'd152;
vramData[13'd1580] = 8'd16;
vramData[13'd1581] = 8'd135;
vramData[13'd1582] = 8'd70;
vramData[13'd1583] = 8'd135;
vramData[13'd1584] = 8'd104;
vramData[13'd1585] = 8'd55;
vramData[13'd1586] = 8'd62;
vramData[13'd1587] = 8'd119;
vramData[13'd1588] = 8'd94;
vramData[13'd1589] = 8'd55;
vramData[13'd1590] = 8'd210;
vramData[13'd1591] = 8'd55;
vramData[13'd1592] = 8'd209;
vramData[13'd1593] = 8'd55;
vramData[13'd1594] = 8'd202;
vramData[13'd1595] = 8'd131;
vramData[13'd1596] = 8'd202;
vramData[13'd1597] = 8'd131;
vramData[13'd1598] = 8'd202;
vramData[13'd1599] = 8'd131;
vramData[13'd1600] = 8'd16;
vramData[13'd1601] = 8'd147;
vramData[13'd1602] = 8'd202;
vramData[13'd1603] = 8'd131;
vramData[13'd1604] = 8'd210;
vramData[13'd1605] = 8'd55;
vramData[13'd1606] = 8'd210;
vramData[13'd1607] = 8'd55;
vramData[13'd1608] = 8'd183;
vramData[13'd1609] = 8'd55;
vramData[13'd1610] = 8'd183;
vramData[13'd1611] = 8'd55;
vramData[13'd1612] = 8'd252;
vramData[13'd1613] = 8'd247;
vramData[13'd1614] = 8'd202;
vramData[13'd1615] = 8'd247;
vramData[13'd1616] = 8'd202;
vramData[13'd1617] = 8'd247;
vramData[13'd1618] = 8'd202;
vramData[13'd1619] = 8'd247;
vramData[13'd1620] = 8'd202;
vramData[13'd1621] = 8'd247;
vramData[13'd1622] = 8'd202;
vramData[13'd1623] = 8'd247;
vramData[13'd1624] = 8'd248;
vramData[13'd1625] = 8'd247;
vramData[13'd1626] = 8'd214;
vramData[13'd1627] = 8'd135;
vramData[13'd1628] = 8'd80;
vramData[13'd1629] = 8'd120;
vramData[13'd1630] = 8'd239;
vramData[13'd1631] = 8'd152;
vramData[13'd1632] = 8'd145;
vramData[13'd1633] = 8'd55;
vramData[13'd1634] = 8'd209;
vramData[13'd1635] = 8'd55;
vramData[13'd1636] = 8'd202;
vramData[13'd1637] = 8'd55;
vramData[13'd1638] = 8'd198;
vramData[13'd1639] = 8'd8;
vramData[13'd1640] = 8'd213;
vramData[13'd1641] = 8'd56;
vramData[13'd1642] = 8'd164;
vramData[13'd1643] = 8'd55;
vramData[13'd1644] = 8'd16;
vramData[13'd1645] = 8'd120;
vramData[13'd1646] = 8'd16;
vramData[13'd1647] = 8'd120;
vramData[13'd1648] = 8'd164;
vramData[13'd1649] = 8'd135;
vramData[13'd1650] = 8'd30;
vramData[13'd1651] = 8'd135;
vramData[13'd1652] = 8'd164;
vramData[13'd1653] = 8'd135;
vramData[13'd1654] = 8'd16;
vramData[13'd1655] = 8'd135;
vramData[13'd1656] = 8'd124;
vramData[13'd1657] = 8'd135;
vramData[13'd1658] = 8'd17;
vramData[13'd1659] = 8'd135;
vramData[13'd1660] = 8'd124;
vramData[13'd1661] = 8'd135;
vramData[13'd1662] = 8'd102;
vramData[13'd1663] = 8'd135;
vramData[13'd1664] = 8'd124;
vramData[13'd1665] = 8'd135;
vramData[13'd1666] = 8'd252;
vramData[13'd1667] = 8'd135;
vramData[13'd1668] = 8'd16;
vramData[13'd1669] = 8'd120;
vramData[13'd1670] = 8'd230;
vramData[13'd1671] = 8'd120;
vramData[13'd1672] = 8'd109;
vramData[13'd1673] = 8'd120;
vramData[13'd1674] = 8'd195;
vramData[13'd1675] = 8'd152;
vramData[13'd1676] = 8'd198;
vramData[13'd1677] = 8'd120;
vramData[13'd1678] = 8'd250;
vramData[13'd1679] = 8'd8;
vramData[13'd1680] = 8'd200;
vramData[13'd1681] = 8'd8;
vramData[13'd1682] = 8'd73;
vramData[13'd1683] = 8'd8;
vramData[13'd1684] = 8'd61;
vramData[13'd1685] = 8'd152;
vramData[13'd1686] = 8'd17;
vramData[13'd1687] = 8'd152;
vramData[13'd1688] = 8'd55;
vramData[13'd1689] = 8'd120;
vramData[13'd1690] = 8'd159;
vramData[13'd1691] = 8'd120;
vramData[13'd1692] = 8'd228;
vramData[13'd1693] = 8'd120;
vramData[13'd1694] = 8'd30;
vramData[13'd1695] = 8'd120;
vramData[13'd1696] = 8'd135;
vramData[13'd1697] = 8'd120;
vramData[13'd1698] = 8'd210;
vramData[13'd1699] = 8'd120;
vramData[13'd1700] = 8'd51;
vramData[13'd1701] = 8'd120;
vramData[13'd1702] = 8'd253;
vramData[13'd1703] = 8'd135;
vramData[13'd1704] = 8'd95;
vramData[13'd1705] = 8'd135;
vramData[13'd1706] = 8'd50;
vramData[13'd1707] = 8'd135;
vramData[13'd1708] = 8'd209;
vramData[13'd1709] = 8'd135;
vramData[13'd1710] = 8'd83;
vramData[13'd1711] = 8'd120;
vramData[13'd1712] = 8'd159;
vramData[13'd1713] = 8'd120;
vramData[13'd1714] = 8'd202;
vramData[13'd1715] = 8'd120;
vramData[13'd1716] = 8'd202;
vramData[13'd1717] = 8'd120;
vramData[13'd1718] = 8'd148;
vramData[13'd1719] = 8'd120;
vramData[13'd1720] = 8'd30;
vramData[13'd1721] = 8'd120;
vramData[13'd1722] = 8'd50;
vramData[13'd1723] = 8'd120;
vramData[13'd1724] = 8'd210;
vramData[13'd1725] = 8'd120;
vramData[13'd1726] = 8'd202;
vramData[13'd1727] = 8'd120;
vramData[13'd1728] = 8'd172;
vramData[13'd1729] = 8'd120;
vramData[13'd1730] = 8'd166;
vramData[13'd1731] = 8'd120;
vramData[13'd1732] = 8'd17;
vramData[13'd1733] = 8'd120;
vramData[13'd1734] = 8'd150;
vramData[13'd1735] = 8'd120;
vramData[13'd1736] = 8'd16;
vramData[13'd1737] = 8'd120;
vramData[13'd1738] = 8'd210;
vramData[13'd1739] = 8'd120;
vramData[13'd1740] = 8'd210;
vramData[13'd1741] = 8'd135;
vramData[13'd1742] = 8'd16;
vramData[13'd1743] = 8'd135;
vramData[13'd1744] = 8'd95;
vramData[13'd1745] = 8'd55;
vramData[13'd1746] = 8'd95;
vramData[13'd1747] = 8'd55;
vramData[13'd1748] = 8'd200;
vramData[13'd1749] = 8'd55;
vramData[13'd1750] = 8'd164;
vramData[13'd1751] = 8'd55;
vramData[13'd1752] = 8'd80;
vramData[13'd1753] = 8'd115;
vramData[13'd1754] = 8'd145;
vramData[13'd1755] = 8'd131;
vramData[13'd1756] = 8'd202;
vramData[13'd1757] = 8'd131;
vramData[13'd1758] = 8'd202;
vramData[13'd1759] = 8'd131;
vramData[13'd1760] = 8'd202;
vramData[13'd1761] = 8'd147;
vramData[13'd1762] = 8'd202;
vramData[13'd1763] = 8'd147;
vramData[13'd1764] = 8'd202;
vramData[13'd1765] = 8'd147;
vramData[13'd1766] = 8'd202;
vramData[13'd1767] = 8'd115;
vramData[13'd1768] = 8'd210;
vramData[13'd1769] = 8'd55;
vramData[13'd1770] = 8'd210;
vramData[13'd1771] = 8'd55;
vramData[13'd1772] = 8'd210;
vramData[13'd1773] = 8'd55;
vramData[13'd1774] = 8'd210;
vramData[13'd1775] = 8'd55;
vramData[13'd1776] = 8'd210;
vramData[13'd1777] = 8'd55;
vramData[13'd1778] = 8'd210;
vramData[13'd1779] = 8'd55;
vramData[13'd1780] = 8'd181;
vramData[13'd1781] = 8'd55;
vramData[13'd1782] = 8'd16;
vramData[13'd1783] = 8'd55;
vramData[13'd1784] = 8'd30;
vramData[13'd1785] = 8'd135;
vramData[13'd1786] = 8'd31;
vramData[13'd1787] = 8'd135;
vramData[13'd1788] = 8'd226;
vramData[13'd1789] = 8'd120;
vramData[13'd1790] = 8'd17;
vramData[13'd1791] = 8'd8;
vramData[13'd1792] = 8'd16;
vramData[13'd1793] = 8'd55;
vramData[13'd1794] = 8'd202;
vramData[13'd1795] = 8'd55;
vramData[13'd1796] = 8'd210;
vramData[13'd1797] = 8'd55;
vramData[13'd1798] = 8'd16;
vramData[13'd1799] = 8'd135;
vramData[13'd1800] = 8'd31;
vramData[13'd1801] = 8'd247;
vramData[13'd1802] = 8'd80;
vramData[13'd1803] = 8'd55;
vramData[13'd1804] = 8'd17;
vramData[13'd1805] = 8'd135;
vramData[13'd1806] = 8'd181;
vramData[13'd1807] = 8'd135;
vramData[13'd1808] = 8'd181;
vramData[13'd1809] = 8'd135;
vramData[13'd1810] = 8'd188;
vramData[13'd1811] = 8'd135;
vramData[13'd1812] = 8'd34;
vramData[13'd1813] = 8'd55;
vramData[13'd1814] = 8'd58;
vramData[13'd1815] = 8'd247;
vramData[13'd1816] = 8'd239;
vramData[13'd1817] = 8'd135;
vramData[13'd1818] = 8'd76;
vramData[13'd1819] = 8'd247;
vramData[13'd1820] = 8'd170;
vramData[13'd1821] = 8'd135;
vramData[13'd1822] = 8'd89;
vramData[13'd1823] = 8'd247;
vramData[13'd1824] = 8'd96;
vramData[13'd1825] = 8'd247;
vramData[13'd1826] = 8'd218;
vramData[13'd1827] = 8'd135;
vramData[13'd1828] = 8'd96;
vramData[13'd1829] = 8'd135;
vramData[13'd1830] = 8'd104;
vramData[13'd1831] = 8'd135;
vramData[13'd1832] = 8'd190;
vramData[13'd1833] = 8'd135;
vramData[13'd1834] = 8'd200;
vramData[13'd1835] = 8'd135;
vramData[13'd1836] = 8'd16;
vramData[13'd1837] = 8'd120;
vramData[13'd1838] = 8'd16;
vramData[13'd1839] = 8'd120;
vramData[13'd1840] = 8'd16;
vramData[13'd1841] = 8'd152;
vramData[13'd1842] = 8'd127;
vramData[13'd1843] = 8'd120;
vramData[13'd1844] = 8'd248;
vramData[13'd1845] = 8'd120;
vramData[13'd1846] = 8'd30;
vramData[13'd1847] = 8'd120;
vramData[13'd1848] = 8'd30;
vramData[13'd1849] = 8'd120;
vramData[13'd1850] = 8'd202;
vramData[13'd1851] = 8'd120;
vramData[13'd1852] = 8'd202;
vramData[13'd1853] = 8'd120;
vramData[13'd1854] = 8'd30;
vramData[13'd1855] = 8'd135;
vramData[13'd1856] = 8'd155;
vramData[13'd1857] = 8'd135;
vramData[13'd1858] = 8'd31;
vramData[13'd1859] = 8'd135;
vramData[13'd1860] = 8'd202;
vramData[13'd1861] = 8'd135;
vramData[13'd1862] = 8'd51;
vramData[13'd1863] = 8'd135;
vramData[13'd1864] = 8'd16;
vramData[13'd1865] = 8'd135;
vramData[13'd1866] = 8'd30;
vramData[13'd1867] = 8'd135;
vramData[13'd1868] = 8'd31;
vramData[13'd1869] = 8'd135;
vramData[13'd1870] = 8'd202;
vramData[13'd1871] = 8'd135;
vramData[13'd1872] = 8'd17;
vramData[13'd1873] = 8'd120;
vramData[13'd1874] = 8'd210;
vramData[13'd1875] = 8'd120;
vramData[13'd1876] = 8'd135;
vramData[13'd1877] = 8'd120;
vramData[13'd1878] = 8'd208;
vramData[13'd1879] = 8'd120;
vramData[13'd1880] = 8'd207;
vramData[13'd1881] = 8'd120;
vramData[13'd1882] = 8'd164;
vramData[13'd1883] = 8'd120;
vramData[13'd1884] = 8'd31;
vramData[13'd1885] = 8'd120;
vramData[13'd1886] = 8'd31;
vramData[13'd1887] = 8'd120;
vramData[13'd1888] = 8'd16;
vramData[13'd1889] = 8'd120;
vramData[13'd1890] = 8'd95;
vramData[13'd1891] = 8'd120;
vramData[13'd1892] = 8'd95;
vramData[13'd1893] = 8'd120;
vramData[13'd1894] = 8'd208;
vramData[13'd1895] = 8'd120;
vramData[13'd1896] = 8'd30;
vramData[13'd1897] = 8'd120;
vramData[13'd1898] = 8'd135;
vramData[13'd1899] = 8'd152;
vramData[13'd1900] = 8'd214;
vramData[13'd1901] = 8'd120;
vramData[13'd1902] = 8'd210;
vramData[13'd1903] = 8'd120;
vramData[13'd1904] = 8'd16;
vramData[13'd1905] = 8'd120;
vramData[13'd1906] = 8'd16;
vramData[13'd1907] = 8'd135;
vramData[13'd1908] = 8'd17;
vramData[13'd1909] = 8'd247;
vramData[13'd1910] = 8'd214;
vramData[13'd1911] = 8'd55;
vramData[13'd1912] = 8'd164;
vramData[13'd1913] = 8'd131;
vramData[13'd1914] = 8'd202;
vramData[13'd1915] = 8'd131;
vramData[13'd1916] = 8'd210;
vramData[13'd1917] = 8'd131;
vramData[13'd1918] = 8'd202;
vramData[13'd1919] = 8'd131;
vramData[13'd1920] = 8'd202;
vramData[13'd1921] = 8'd147;
vramData[13'd1922] = 8'd202;
vramData[13'd1923] = 8'd147;
vramData[13'd1924] = 8'd202;
vramData[13'd1925] = 8'd147;
vramData[13'd1926] = 8'd202;
vramData[13'd1927] = 8'd147;
vramData[13'd1928] = 8'd202;
vramData[13'd1929] = 8'd147;
vramData[13'd1930] = 8'd202;
vramData[13'd1931] = 8'd147;
vramData[13'd1932] = 8'd202;
vramData[13'd1933] = 8'd147;
vramData[13'd1934] = 8'd202;
vramData[13'd1935] = 8'd147;
vramData[13'd1936] = 8'd202;
vramData[13'd1937] = 8'd147;
vramData[13'd1938] = 8'd202;
vramData[13'd1939] = 8'd147;
vramData[13'd1940] = 8'd210;
vramData[13'd1941] = 8'd135;
vramData[13'd1942] = 8'd164;
vramData[13'd1943] = 8'd120;
vramData[13'd1944] = 8'd16;
vramData[13'd1945] = 8'd135;
vramData[13'd1946] = 8'd209;
vramData[13'd1947] = 8'd135;
vramData[13'd1948] = 8'd16;
vramData[13'd1949] = 8'd120;
vramData[13'd1950] = 8'd200;
vramData[13'd1951] = 8'd8;
vramData[13'd1952] = 8'd30;
vramData[13'd1953] = 8'd8;
vramData[13'd1954] = 8'd202;
vramData[13'd1955] = 8'd56;
vramData[13'd1956] = 8'd202;
vramData[13'd1957] = 8'd115;
vramData[13'd1958] = 8'd210;
vramData[13'd1959] = 8'd55;
vramData[13'd1960] = 8'd210;
vramData[13'd1961] = 8'd55;
vramData[13'd1962] = 8'd198;
vramData[13'd1963] = 8'd135;
vramData[13'd1964] = 8'd214;
vramData[13'd1965] = 8'd135;
vramData[13'd1966] = 8'd145;
vramData[13'd1967] = 8'd135;
vramData[13'd1968] = 8'd135;
vramData[13'd1969] = 8'd135;
vramData[13'd1970] = 8'd104;
vramData[13'd1971] = 8'd135;
vramData[13'd1972] = 8'd7;
vramData[13'd1973] = 8'd247;
vramData[13'd1974] = 8'd28;
vramData[13'd1975] = 8'd135;
vramData[13'd1976] = 8'd164;
vramData[13'd1977] = 8'd247;
vramData[13'd1978] = 8'd109;
vramData[13'd1979] = 8'd247;
vramData[13'd1980] = 8'd9;
vramData[13'd1981] = 8'd247;
vramData[13'd1982] = 8'd39;
vramData[13'd1983] = 8'd247;
vramData[13'd1984] = 8'd24;
vramData[13'd1985] = 8'd103;
vramData[13'd1986] = 8'd16;
vramData[13'd1987] = 8'd247;
vramData[13'd1988] = 8'd17;
vramData[13'd1989] = 8'd247;
vramData[13'd1990] = 8'd17;
vramData[13'd1991] = 8'd247;
vramData[13'd1992] = 8'd95;
vramData[13'd1993] = 8'd247;
vramData[13'd1994] = 8'd39;
vramData[13'd1995] = 8'd135;
vramData[13'd1996] = 8'd16;
vramData[13'd1997] = 8'd120;
vramData[13'd1998] = 8'd80;
vramData[13'd1999] = 8'd120;
vramData[13'd2000] = 8'd94;
vramData[13'd2001] = 8'd152;
vramData[13'd2002] = 8'd214;
vramData[13'd2003] = 8'd8;
vramData[13'd2004] = 8'd31;
vramData[13'd2005] = 8'd8;
vramData[13'd2006] = 8'd202;
vramData[13'd2007] = 8'd8;
vramData[13'd2008] = 8'd95;
vramData[13'd2009] = 8'd56;
vramData[13'd2010] = 8'd214;
vramData[13'd2011] = 8'd152;
vramData[13'd2012] = 8'd95;
vramData[13'd2013] = 8'd56;
vramData[13'd2014] = 8'd95;
vramData[13'd2015] = 8'd56;
vramData[13'd2016] = 8'd95;
vramData[13'd2017] = 8'd56;
vramData[13'd2018] = 8'd126;
vramData[13'd2019] = 8'd120;
vramData[13'd2020] = 8'd200;
vramData[13'd2021] = 8'd120;
vramData[13'd2022] = 8'd30;
vramData[13'd2023] = 8'd120;
vramData[13'd2024] = 8'd83;
vramData[13'd2025] = 8'd120;
vramData[13'd2026] = 8'd239;
vramData[13'd2027] = 8'd135;
vramData[13'd2028] = 8'd167;
vramData[13'd2029] = 8'd135;
vramData[13'd2030] = 8'd166;
vramData[13'd2031] = 8'd135;
vramData[13'd2032] = 8'd226;
vramData[13'd2033] = 8'd135;
vramData[13'd2034] = 8'd240;
vramData[13'd2035] = 8'd120;
vramData[13'd2036] = 8'd17;
vramData[13'd2037] = 8'd120;
vramData[13'd2038] = 8'd80;
vramData[13'd2039] = 8'd120;
vramData[13'd2040] = 8'd181;
vramData[13'd2041] = 8'd120;
vramData[13'd2042] = 8'd37;
vramData[13'd2043] = 8'd120;
vramData[13'd2044] = 8'd16;
vramData[13'd2045] = 8'd120;
vramData[13'd2046] = 8'd31;
vramData[13'd2047] = 8'd120;
vramData[13'd2048] = 8'd83;
vramData[13'd2049] = 8'd120;
vramData[13'd2050] = 8'd210;
vramData[13'd2051] = 8'd120;
vramData[13'd2052] = 8'd17;
vramData[13'd2053] = 8'd120;
vramData[13'd2054] = 8'd202;
vramData[13'd2055] = 8'd120;
vramData[13'd2056] = 8'd31;
vramData[13'd2057] = 8'd120;
vramData[13'd2058] = 8'd70;
vramData[13'd2059] = 8'd120;
vramData[13'd2060] = 8'd208;
vramData[13'd2061] = 8'd120;
vramData[13'd2062] = 8'd210;
vramData[13'd2063] = 8'd120;
vramData[13'd2064] = 8'd223;
vramData[13'd2065] = 8'd135;
vramData[13'd2066] = 8'd214;
vramData[13'd2067] = 8'd55;
vramData[13'd2068] = 8'd80;
vramData[13'd2069] = 8'd120;
vramData[13'd2070] = 8'd202;
vramData[13'd2071] = 8'd56;
vramData[13'd2072] = 8'd202;
vramData[13'd2073] = 8'd56;
vramData[13'd2074] = 8'd202;
vramData[13'd2075] = 8'd56;
vramData[13'd2076] = 8'd202;
vramData[13'd2077] = 8'd56;
vramData[13'd2078] = 8'd202;
vramData[13'd2079] = 8'd56;
vramData[13'd2080] = 8'd202;
vramData[13'd2081] = 8'd24;
vramData[13'd2082] = 8'd202;
vramData[13'd2083] = 8'd24;
vramData[13'd2084] = 8'd202;
vramData[13'd2085] = 8'd24;
vramData[13'd2086] = 8'd202;
vramData[13'd2087] = 8'd24;
vramData[13'd2088] = 8'd202;
vramData[13'd2089] = 8'd24;
vramData[13'd2090] = 8'd210;
vramData[13'd2091] = 8'd8;
vramData[13'd2092] = 8'd210;
vramData[13'd2093] = 8'd8;
vramData[13'd2094] = 8'd16;
vramData[13'd2095] = 8'd8;
vramData[13'd2096] = 8'd202;
vramData[13'd2097] = 8'd56;
vramData[13'd2098] = 8'd202;
vramData[13'd2099] = 8'd56;
vramData[13'd2100] = 8'd80;
vramData[13'd2101] = 8'd152;
vramData[13'd2102] = 8'd202;
vramData[13'd2103] = 8'd152;
vramData[13'd2104] = 8'd202;
vramData[13'd2105] = 8'd152;
vramData[13'd2106] = 8'd51;
vramData[13'd2107] = 8'd120;
vramData[13'd2108] = 8'd210;
vramData[13'd2109] = 8'd135;
vramData[13'd2110] = 8'd208;
vramData[13'd2111] = 8'd135;
vramData[13'd2112] = 8'd202;
vramData[13'd2113] = 8'd135;
vramData[13'd2114] = 8'd220;
vramData[13'd2115] = 8'd120;
vramData[13'd2116] = 8'd210;
vramData[13'd2117] = 8'd120;
vramData[13'd2118] = 8'd210;
vramData[13'd2119] = 8'd120;
vramData[13'd2120] = 8'd31;
vramData[13'd2121] = 8'd135;
vramData[13'd2122] = 8'd31;
vramData[13'd2123] = 8'd135;
vramData[13'd2124] = 8'd220;
vramData[13'd2125] = 8'd120;
vramData[13'd2126] = 8'd253;
vramData[13'd2127] = 8'd135;
vramData[13'd2128] = 8'd205;
vramData[13'd2129] = 8'd135;
vramData[13'd2130] = 8'd95;
vramData[13'd2131] = 8'd247;
vramData[13'd2132] = 8'd89;
vramData[13'd2133] = 8'd247;
vramData[13'd2134] = 8'd202;
vramData[13'd2135] = 8'd247;
vramData[13'd2136] = 8'd19;
vramData[13'd2137] = 8'd247;
vramData[13'd2138] = 8'd89;
vramData[13'd2139] = 8'd247;
vramData[13'd2140] = 8'd93;
vramData[13'd2141] = 8'd247;
vramData[13'd2142] = 8'd245;
vramData[13'd2143] = 8'd247;
vramData[13'd2144] = 8'd200;
vramData[13'd2145] = 8'd247;
vramData[13'd2146] = 8'd129;
vramData[13'd2147] = 8'd247;
vramData[13'd2148] = 8'd30;
vramData[13'd2149] = 8'd247;
vramData[13'd2150] = 8'd86;
vramData[13'd2151] = 8'd247;
vramData[13'd2152] = 8'd33;
vramData[13'd2153] = 8'd87;
vramData[13'd2154] = 8'd31;
vramData[13'd2155] = 8'd135;
vramData[13'd2156] = 8'd171;
vramData[13'd2157] = 8'd120;
vramData[13'd2158] = 8'd95;
vramData[13'd2159] = 8'd8;
vramData[13'd2160] = 8'd214;
vramData[13'd2161] = 8'd8;
vramData[13'd2162] = 8'd16;
vramData[13'd2163] = 8'd8;
vramData[13'd2164] = 8'd80;
vramData[13'd2165] = 8'd135;
vramData[13'd2166] = 8'd202;
vramData[13'd2167] = 8'd55;
vramData[13'd2168] = 8'd202;
vramData[13'd2169] = 8'd55;
vramData[13'd2170] = 8'd31;
vramData[13'd2171] = 8'd115;
vramData[13'd2172] = 8'd16;
vramData[13'd2173] = 8'd120;
vramData[13'd2174] = 8'd31;
vramData[13'd2175] = 8'd8;
vramData[13'd2176] = 8'd198;
vramData[13'd2177] = 8'd120;
vramData[13'd2178] = 8'd16;
vramData[13'd2179] = 8'd55;
vramData[13'd2180] = 8'd209;
vramData[13'd2181] = 8'd55;
vramData[13'd2182] = 8'd183;
vramData[13'd2183] = 8'd120;
vramData[13'd2184] = 8'd230;
vramData[13'd2185] = 8'd152;
vramData[13'd2186] = 8'd200;
vramData[13'd2187] = 8'd120;
vramData[13'd2188] = 8'd83;
vramData[13'd2189] = 8'd135;
vramData[13'd2190] = 8'd16;
vramData[13'd2191] = 8'd135;
vramData[13'd2192] = 8'd50;
vramData[13'd2193] = 8'd135;
vramData[13'd2194] = 8'd80;
vramData[13'd2195] = 8'd135;
vramData[13'd2196] = 8'd17;
vramData[13'd2197] = 8'd120;
vramData[13'd2198] = 8'd198;
vramData[13'd2199] = 8'd120;
vramData[13'd2200] = 8'd210;
vramData[13'd2201] = 8'd120;
vramData[13'd2202] = 8'd80;
vramData[13'd2203] = 8'd120;
vramData[13'd2204] = 8'd51;
vramData[13'd2205] = 8'd120;
vramData[13'd2206] = 8'd156;
vramData[13'd2207] = 8'd120;
vramData[13'd2208] = 8'd51;
vramData[13'd2209] = 8'd120;
vramData[13'd2210] = 8'd17;
vramData[13'd2211] = 8'd120;
vramData[13'd2212] = 8'd214;
vramData[13'd2213] = 8'd120;
vramData[13'd2214] = 8'd17;
vramData[13'd2215] = 8'd120;
vramData[13'd2216] = 8'd202;
vramData[13'd2217] = 8'd120;
vramData[13'd2218] = 8'd171;
vramData[13'd2219] = 8'd120;
vramData[13'd2220] = 8'd214;
vramData[13'd2221] = 8'd120;
vramData[13'd2222] = 8'd226;
vramData[13'd2223] = 8'd135;
vramData[13'd2224] = 8'd226;
vramData[13'd2225] = 8'd247;
vramData[13'd2226] = 8'd198;
vramData[13'd2227] = 8'd55;
vramData[13'd2228] = 8'd16;
vramData[13'd2229] = 8'd147;
vramData[13'd2230] = 8'd202;
vramData[13'd2231] = 8'd19;
vramData[13'd2232] = 8'd202;
vramData[13'd2233] = 8'd19;
vramData[13'd2234] = 8'd202;
vramData[13'd2235] = 8'd19;
vramData[13'd2236] = 8'd202;
vramData[13'd2237] = 8'd19;
vramData[13'd2238] = 8'd202;
vramData[13'd2239] = 8'd19;
vramData[13'd2240] = 8'd210;
vramData[13'd2241] = 8'd115;
vramData[13'd2242] = 8'd202;
vramData[13'd2243] = 8'd131;
vramData[13'd2244] = 8'd202;
vramData[13'd2245] = 8'd131;
vramData[13'd2246] = 8'd210;
vramData[13'd2247] = 8'd56;
vramData[13'd2248] = 8'd164;
vramData[13'd2249] = 8'd24;
vramData[13'd2250] = 8'd202;
vramData[13'd2251] = 8'd24;
vramData[13'd2252] = 8'd80;
vramData[13'd2253] = 8'd8;
vramData[13'd2254] = 8'd95;
vramData[13'd2255] = 8'd8;
vramData[13'd2256] = 8'd202;
vramData[13'd2257] = 8'd152;
vramData[13'd2258] = 8'd202;
vramData[13'd2259] = 8'd152;
vramData[13'd2260] = 8'd202;
vramData[13'd2261] = 8'd152;
vramData[13'd2262] = 8'd135;
vramData[13'd2263] = 8'd152;
vramData[13'd2264] = 8'd202;
vramData[13'd2265] = 8'd152;
vramData[13'd2266] = 8'd109;
vramData[13'd2267] = 8'd152;
vramData[13'd2268] = 8'd166;
vramData[13'd2269] = 8'd120;
vramData[13'd2270] = 8'd16;
vramData[13'd2271] = 8'd135;
vramData[13'd2272] = 8'd135;
vramData[13'd2273] = 8'd135;
vramData[13'd2274] = 8'd16;
vramData[13'd2275] = 8'd135;
vramData[13'd2276] = 8'd31;
vramData[13'd2277] = 8'd55;
vramData[13'd2278] = 8'd80;
vramData[13'd2279] = 8'd55;
vramData[13'd2280] = 8'd183;
vramData[13'd2281] = 8'd247;
vramData[13'd2282] = 8'd51;
vramData[13'd2283] = 8'd247;
vramData[13'd2284] = 8'd226;
vramData[13'd2285] = 8'd247;
vramData[13'd2286] = 8'd70;
vramData[13'd2287] = 8'd247;
vramData[13'd2288] = 8'd52;
vramData[13'd2289] = 8'd247;
vramData[13'd2290] = 8'd167;
vramData[13'd2291] = 8'd247;
vramData[13'd2292] = 8'd107;
vramData[13'd2293] = 8'd247;
vramData[13'd2294] = 8'd119;
vramData[13'd2295] = 8'd247;
vramData[13'd2296] = 8'd190;
vramData[13'd2297] = 8'd247;
vramData[13'd2298] = 8'd16;
vramData[13'd2299] = 8'd247;
vramData[13'd2300] = 8'd16;
vramData[13'd2301] = 8'd247;
vramData[13'd2302] = 8'd30;
vramData[13'd2303] = 8'd247;
vramData[13'd2304] = 8'd156;
vramData[13'd2305] = 8'd247;
vramData[13'd2306] = 8'd202;
vramData[13'd2307] = 8'd247;
vramData[13'd2308] = 8'd75;
vramData[13'd2309] = 8'd247;
vramData[13'd2310] = 8'd24;
vramData[13'd2311] = 8'd87;
vramData[13'd2312] = 8'd218;
vramData[13'd2313] = 8'd247;
vramData[13'd2314] = 8'd226;
vramData[13'd2315] = 8'd120;
vramData[13'd2316] = 8'd210;
vramData[13'd2317] = 8'd8;
vramData[13'd2318] = 8'd37;
vramData[13'd2319] = 8'd128;
vramData[13'd2320] = 8'd164;
vramData[13'd2321] = 8'd8;
vramData[13'd2322] = 8'd221;
vramData[13'd2323] = 8'd135;
vramData[13'd2324] = 8'd209;
vramData[13'd2325] = 8'd183;
vramData[13'd2326] = 8'd16;
vramData[13'd2327] = 8'd183;
vramData[13'd2328] = 8'd17;
vramData[13'd2329] = 8'd183;
vramData[13'd2330] = 8'd16;
vramData[13'd2331] = 8'd183;
vramData[13'd2332] = 8'd16;
vramData[13'd2333] = 8'd8;
vramData[13'd2334] = 8'd16;
vramData[13'd2335] = 8'd8;
vramData[13'd2336] = 8'd80;
vramData[13'd2337] = 8'd135;
vramData[13'd2338] = 8'd80;
vramData[13'd2339] = 8'd183;
vramData[13'd2340] = 8'd16;
vramData[13'd2341] = 8'd183;
vramData[13'd2342] = 8'd31;
vramData[13'd2343] = 8'd247;
vramData[13'd2344] = 8'd200;
vramData[13'd2345] = 8'd55;
vramData[13'd2346] = 8'd16;
vramData[13'd2347] = 8'd120;
vramData[13'd2348] = 8'd17;
vramData[13'd2349] = 8'd120;
vramData[13'd2350] = 8'd16;
vramData[13'd2351] = 8'd135;
vramData[13'd2352] = 8'd164;
vramData[13'd2353] = 8'd135;
vramData[13'd2354] = 8'd83;
vramData[13'd2355] = 8'd120;
vramData[13'd2356] = 8'd209;
vramData[13'd2357] = 8'd120;
vramData[13'd2358] = 8'd37;
vramData[13'd2359] = 8'd135;
vramData[13'd2360] = 8'd202;
vramData[13'd2361] = 8'd135;
vramData[13'd2362] = 8'd31;
vramData[13'd2363] = 8'd120;
vramData[13'd2364] = 8'd197;
vramData[13'd2365] = 8'd120;
vramData[13'd2366] = 8'd9;
vramData[13'd2367] = 8'd120;
vramData[13'd2368] = 8'd31;
vramData[13'd2369] = 8'd135;
vramData[13'd2370] = 8'd31;
vramData[13'd2371] = 8'd135;
vramData[13'd2372] = 8'd61;
vramData[13'd2373] = 8'd135;
vramData[13'd2374] = 8'd200;
vramData[13'd2375] = 8'd135;
vramData[13'd2376] = 8'd202;
vramData[13'd2377] = 8'd135;
vramData[13'd2378] = 8'd202;
vramData[13'd2379] = 8'd135;
vramData[13'd2380] = 8'd253;
vramData[13'd2381] = 8'd135;
vramData[13'd2382] = 8'd75;
vramData[13'd2383] = 8'd119;
vramData[13'd2384] = 8'd16;
vramData[13'd2385] = 8'd87;
vramData[13'd2386] = 8'd198;
vramData[13'd2387] = 8'd55;
vramData[13'd2388] = 8'd210;
vramData[13'd2389] = 8'd147;
vramData[13'd2390] = 8'd16;
vramData[13'd2391] = 8'd147;
vramData[13'd2392] = 8'd210;
vramData[13'd2393] = 8'd147;
vramData[13'd2394] = 8'd210;
vramData[13'd2395] = 8'd147;
vramData[13'd2396] = 8'd210;
vramData[13'd2397] = 8'd147;
vramData[13'd2398] = 8'd210;
vramData[13'd2399] = 8'd147;
vramData[13'd2400] = 8'd210;
vramData[13'd2401] = 8'd147;
vramData[13'd2402] = 8'd210;
vramData[13'd2403] = 8'd147;
vramData[13'd2404] = 8'd210;
vramData[13'd2405] = 8'd147;
vramData[13'd2406] = 8'd202;
vramData[13'd2407] = 8'd131;
vramData[13'd2408] = 8'd16;
vramData[13'd2409] = 8'd56;
vramData[13'd2410] = 8'd145;
vramData[13'd2411] = 8'd24;
vramData[13'd2412] = 8'd202;
vramData[13'd2413] = 8'd8;
vramData[13'd2414] = 8'd31;
vramData[13'd2415] = 8'd8;
vramData[13'd2416] = 8'd16;
vramData[13'd2417] = 8'd8;
vramData[13'd2418] = 8'd214;
vramData[13'd2419] = 8'd152;
vramData[13'd2420] = 8'd181;
vramData[13'd2421] = 8'd152;
vramData[13'd2422] = 8'd85;
vramData[13'd2423] = 8'd152;
vramData[13'd2424] = 8'd210;
vramData[13'd2425] = 8'd152;
vramData[13'd2426] = 8'd214;
vramData[13'd2427] = 8'd120;
vramData[13'd2428] = 8'd80;
vramData[13'd2429] = 8'd135;
vramData[13'd2430] = 8'd202;
vramData[13'd2431] = 8'd135;
vramData[13'd2432] = 8'd31;
vramData[13'd2433] = 8'd55;
vramData[13'd2434] = 8'd202;
vramData[13'd2435] = 8'd55;
vramData[13'd2436] = 8'd248;
vramData[13'd2437] = 8'd55;
vramData[13'd2438] = 8'd37;
vramData[13'd2439] = 8'd247;
vramData[13'd2440] = 8'd230;
vramData[13'd2441] = 8'd247;
vramData[13'd2442] = 8'd241;
vramData[13'd2443] = 8'd247;
vramData[13'd2444] = 8'd210;
vramData[13'd2445] = 8'd247;
vramData[13'd2446] = 8'd240;
vramData[13'd2447] = 8'd247;
vramData[13'd2448] = 8'd171;
vramData[13'd2449] = 8'd247;
vramData[13'd2450] = 8'd31;
vramData[13'd2451] = 8'd247;
vramData[13'd2452] = 8'd86;
vramData[13'd2453] = 8'd247;
vramData[13'd2454] = 8'd106;
vramData[13'd2455] = 8'd247;
vramData[13'd2456] = 8'd181;
vramData[13'd2457] = 8'd247;
vramData[13'd2458] = 8'd7;
vramData[13'd2459] = 8'd247;
vramData[13'd2460] = 8'd239;
vramData[13'd2461] = 8'd247;
vramData[13'd2462] = 8'd252;
vramData[13'd2463] = 8'd247;
vramData[13'd2464] = 8'd198;
vramData[13'd2465] = 8'd87;
vramData[13'd2466] = 8'd31;
vramData[13'd2467] = 8'd135;
vramData[13'd2468] = 8'd240;
vramData[13'd2469] = 8'd247;
vramData[13'd2470] = 8'd218;
vramData[13'd2471] = 8'd247;
vramData[13'd2472] = 8'd188;
vramData[13'd2473] = 8'd247;
vramData[13'd2474] = 8'd202;
vramData[13'd2475] = 8'd135;
vramData[13'd2476] = 8'd200;
vramData[13'd2477] = 8'd8;
vramData[13'd2478] = 8'd16;
vramData[13'd2479] = 8'd128;
vramData[13'd2480] = 8'd17;
vramData[13'd2481] = 8'd128;
vramData[13'd2482] = 8'd200;
vramData[13'd2483] = 8'd120;
vramData[13'd2484] = 8'd202;
vramData[13'd2485] = 8'd183;
vramData[13'd2486] = 8'd164;
vramData[13'd2487] = 8'd183;
vramData[13'd2488] = 8'd209;
vramData[13'd2489] = 8'd183;
vramData[13'd2490] = 8'd181;
vramData[13'd2491] = 8'd183;
vramData[13'd2492] = 8'd223;
vramData[13'd2493] = 8'd135;
vramData[13'd2494] = 8'd70;
vramData[13'd2495] = 8'd135;
vramData[13'd2496] = 8'd37;
vramData[13'd2497] = 8'd247;
vramData[13'd2498] = 8'd30;
vramData[13'd2499] = 8'd183;
vramData[13'd2500] = 8'd210;
vramData[13'd2501] = 8'd183;
vramData[13'd2502] = 8'd16;
vramData[13'd2503] = 8'd183;
vramData[13'd2504] = 8'd220;
vramData[13'd2505] = 8'd135;
vramData[13'd2506] = 8'd76;
vramData[13'd2507] = 8'd152;
vramData[13'd2508] = 8'd67;
vramData[13'd2509] = 8'd135;
vramData[13'd2510] = 8'd17;
vramData[13'd2511] = 8'd135;
vramData[13'd2512] = 8'd171;
vramData[13'd2513] = 8'd120;
vramData[13'd2514] = 8'd202;
vramData[13'd2515] = 8'd120;
vramData[13'd2516] = 8'd117;
vramData[13'd2517] = 8'd120;
vramData[13'd2518] = 8'd37;
vramData[13'd2519] = 8'd120;
vramData[13'd2520] = 8'd30;
vramData[13'd2521] = 8'd135;
vramData[13'd2522] = 8'd240;
vramData[13'd2523] = 8'd120;
vramData[13'd2524] = 8'd156;
vramData[13'd2525] = 8'd135;
vramData[13'd2526] = 8'd240;
vramData[13'd2527] = 8'd135;
vramData[13'd2528] = 8'd240;
vramData[13'd2529] = 8'd135;
vramData[13'd2530] = 8'd30;
vramData[13'd2531] = 8'd135;
vramData[13'd2532] = 8'd17;
vramData[13'd2533] = 8'd135;
vramData[13'd2534] = 8'd46;
vramData[13'd2535] = 8'd135;
vramData[13'd2536] = 8'd126;
vramData[13'd2537] = 8'd135;
vramData[13'd2538] = 8'd135;
vramData[13'd2539] = 8'd55;
vramData[13'd2540] = 8'd16;
vramData[13'd2541] = 8'd55;
vramData[13'd2542] = 8'd71;
vramData[13'd2543] = 8'd119;
vramData[13'd2544] = 8'd117;
vramData[13'd2545] = 8'd247;
vramData[13'd2546] = 8'd16;
vramData[13'd2547] = 8'd247;
vramData[13'd2548] = 8'd16;
vramData[13'd2549] = 8'd115;
vramData[13'd2550] = 8'd145;
vramData[13'd2551] = 8'd179;
vramData[13'd2552] = 8'd145;
vramData[13'd2553] = 8'd179;
vramData[13'd2554] = 8'd145;
vramData[13'd2555] = 8'd179;
vramData[13'd2556] = 8'd145;
vramData[13'd2557] = 8'd179;
vramData[13'd2558] = 8'd16;
vramData[13'd2559] = 8'd179;
vramData[13'd2560] = 8'd210;
vramData[13'd2561] = 8'd147;
vramData[13'd2562] = 8'd181;
vramData[13'd2563] = 8'd147;
vramData[13'd2564] = 8'd202;
vramData[13'd2565] = 8'd147;
vramData[13'd2566] = 8'd164;
vramData[13'd2567] = 8'd147;
vramData[13'd2568] = 8'd202;
vramData[13'd2569] = 8'd131;
vramData[13'd2570] = 8'd202;
vramData[13'd2571] = 8'd131;
vramData[13'd2572] = 8'd145;
vramData[13'd2573] = 8'd24;
vramData[13'd2574] = 8'd214;
vramData[13'd2575] = 8'd152;
vramData[13'd2576] = 8'd70;
vramData[13'd2577] = 8'd135;
vramData[13'd2578] = 8'd200;
vramData[13'd2579] = 8'd135;
vramData[13'd2580] = 8'd16;
vramData[13'd2581] = 8'd120;
vramData[13'd2582] = 8'd210;
vramData[13'd2583] = 8'd120;
vramData[13'd2584] = 8'd210;
vramData[13'd2585] = 8'd120;
vramData[13'd2586] = 8'd16;
vramData[13'd2587] = 8'd135;
vramData[13'd2588] = 8'd164;
vramData[13'd2589] = 8'd55;
vramData[13'd2590] = 8'd30;
vramData[13'd2591] = 8'd55;
vramData[13'd2592] = 8'd214;
vramData[13'd2593] = 8'd247;
vramData[13'd2594] = 8'd9;
vramData[13'd2595] = 8'd247;
vramData[13'd2596] = 8'd107;
vramData[13'd2597] = 8'd247;
vramData[13'd2598] = 8'd241;
vramData[13'd2599] = 8'd247;
vramData[13'd2600] = 8'd31;
vramData[13'd2601] = 8'd247;
vramData[13'd2602] = 8'd157;
vramData[13'd2603] = 8'd247;
vramData[13'd2604] = 8'd83;
vramData[13'd2605] = 8'd247;
vramData[13'd2606] = 8'd83;
vramData[13'd2607] = 8'd247;
vramData[13'd2608] = 8'd37;
vramData[13'd2609] = 8'd247;
vramData[13'd2610] = 8'd109;
vramData[13'd2611] = 8'd247;
vramData[13'd2612] = 8'd108;
vramData[13'd2613] = 8'd247;
vramData[13'd2614] = 8'd252;
vramData[13'd2615] = 8'd247;
vramData[13'd2616] = 8'd159;
vramData[13'd2617] = 8'd247;
vramData[13'd2618] = 8'd86;
vramData[13'd2619] = 8'd247;
vramData[13'd2620] = 8'd95;
vramData[13'd2621] = 8'd135;
vramData[13'd2622] = 8'd52;
vramData[13'd2623] = 8'd135;
vramData[13'd2624] = 8'd52;
vramData[13'd2625] = 8'd135;
vramData[13'd2626] = 8'd16;
vramData[13'd2627] = 8'd135;
vramData[13'd2628] = 8'd127;
vramData[13'd2629] = 8'd135;
vramData[13'd2630] = 8'd28;
vramData[13'd2631] = 8'd135;
vramData[13'd2632] = 8'd183;
vramData[13'd2633] = 8'd87;
vramData[13'd2634] = 8'd16;
vramData[13'd2635] = 8'd87;
vramData[13'd2636] = 8'd46;
vramData[13'd2637] = 8'd135;
vramData[13'd2638] = 8'd200;
vramData[13'd2639] = 8'd135;
vramData[13'd2640] = 8'd183;
vramData[13'd2641] = 8'd120;
vramData[13'd2642] = 8'd166;
vramData[13'd2643] = 8'd8;
vramData[13'd2644] = 8'd202;
vramData[13'd2645] = 8'd56;
vramData[13'd2646] = 8'd223;
vramData[13'd2647] = 8'd120;
vramData[13'd2648] = 8'd145;
vramData[13'd2649] = 8'd183;
vramData[13'd2650] = 8'd145;
vramData[13'd2651] = 8'd183;
vramData[13'd2652] = 8'd210;
vramData[13'd2653] = 8'd55;
vramData[13'd2654] = 8'd210;
vramData[13'd2655] = 8'd55;
vramData[13'd2656] = 8'd210;
vramData[13'd2657] = 8'd55;
vramData[13'd2658] = 8'd202;
vramData[13'd2659] = 8'd115;
vramData[13'd2660] = 8'd80;
vramData[13'd2661] = 8'd56;
vramData[13'd2662] = 8'd95;
vramData[13'd2663] = 8'd120;
vramData[13'd2664] = 8'd214;
vramData[13'd2665] = 8'd120;
vramData[13'd2666] = 8'd107;
vramData[13'd2667] = 8'd135;
vramData[13'd2668] = 8'd164;
vramData[13'd2669] = 8'd135;
vramData[13'd2670] = 8'd67;
vramData[13'd2671] = 8'd135;
vramData[13'd2672] = 8'd18;
vramData[13'd2673] = 8'd135;
vramData[13'd2674] = 8'd210;
vramData[13'd2675] = 8'd135;
vramData[13'd2676] = 8'd210;
vramData[13'd2677] = 8'd120;
vramData[13'd2678] = 8'd210;
vramData[13'd2679] = 8'd120;
vramData[13'd2680] = 8'd30;
vramData[13'd2681] = 8'd120;
vramData[13'd2682] = 8'd90;
vramData[13'd2683] = 8'd120;
vramData[13'd2684] = 8'd101;
vramData[13'd2685] = 8'd120;
vramData[13'd2686] = 8'd240;
vramData[13'd2687] = 8'd135;
vramData[13'd2688] = 8'd240;
vramData[13'd2689] = 8'd135;
vramData[13'd2690] = 8'd240;
vramData[13'd2691] = 8'd135;
vramData[13'd2692] = 8'd28;
vramData[13'd2693] = 8'd135;
vramData[13'd2694] = 8'd226;
vramData[13'd2695] = 8'd135;
vramData[13'd2696] = 8'd51;
vramData[13'd2697] = 8'd55;
vramData[13'd2698] = 8'd31;
vramData[13'd2699] = 8'd55;
vramData[13'd2700] = 8'd92;
vramData[13'd2701] = 8'd55;
vramData[13'd2702] = 8'd95;
vramData[13'd2703] = 8'd247;
vramData[13'd2704] = 8'd192;
vramData[13'd2705] = 8'd119;
vramData[13'd2706] = 8'd30;
vramData[13'd2707] = 8'd247;
vramData[13'd2708] = 8'd222;
vramData[13'd2709] = 8'd135;
vramData[13'd2710] = 8'd202;
vramData[13'd2711] = 8'd56;
vramData[13'd2712] = 8'd223;
vramData[13'd2713] = 8'd56;
vramData[13'd2714] = 8'd220;
vramData[13'd2715] = 8'd131;
vramData[13'd2716] = 8'd220;
vramData[13'd2717] = 8'd131;
vramData[13'd2718] = 8'd220;
vramData[13'd2719] = 8'd131;
vramData[13'd2720] = 8'd202;
vramData[13'd2721] = 8'd147;
vramData[13'd2722] = 8'd202;
vramData[13'd2723] = 8'd147;
vramData[13'd2724] = 8'd181;
vramData[13'd2725] = 8'd147;
vramData[13'd2726] = 8'd210;
vramData[13'd2727] = 8'd147;
vramData[13'd2728] = 8'd210;
vramData[13'd2729] = 8'd147;
vramData[13'd2730] = 8'd202;
vramData[13'd2731] = 8'd131;
vramData[13'd2732] = 8'd210;
vramData[13'd2733] = 8'd56;
vramData[13'd2734] = 8'd70;
vramData[13'd2735] = 8'd55;
vramData[13'd2736] = 8'd183;
vramData[13'd2737] = 8'd247;
vramData[13'd2738] = 8'd95;
vramData[13'd2739] = 8'd247;
vramData[13'd2740] = 8'd200;
vramData[13'd2741] = 8'd135;
vramData[13'd2742] = 8'd202;
vramData[13'd2743] = 8'd135;
vramData[13'd2744] = 8'd210;
vramData[13'd2745] = 8'd135;
vramData[13'd2746] = 8'd210;
vramData[13'd2747] = 8'd55;
vramData[13'd2748] = 8'd230;
vramData[13'd2749] = 8'd55;
vramData[13'd2750] = 8'd95;
vramData[13'd2751] = 8'd135;
vramData[13'd2752] = 8'd210;
vramData[13'd2753] = 8'd55;
vramData[13'd2754] = 8'd28;
vramData[13'd2755] = 8'd55;
vramData[13'd2756] = 8'd228;
vramData[13'd2757] = 8'd55;
vramData[13'd2758] = 8'd253;
vramData[13'd2759] = 8'd247;
vramData[13'd2760] = 8'd162;
vramData[13'd2761] = 8'd247;
vramData[13'd2762] = 8'd197;
vramData[13'd2763] = 8'd247;
vramData[13'd2764] = 8'd202;
vramData[13'd2765] = 8'd247;
vramData[13'd2766] = 8'd239;
vramData[13'd2767] = 8'd247;
vramData[13'd2768] = 8'd202;
vramData[13'd2769] = 8'd247;
vramData[13'd2770] = 8'd252;
vramData[13'd2771] = 8'd247;
vramData[13'd2772] = 8'd253;
vramData[13'd2773] = 8'd247;
vramData[13'd2774] = 8'd102;
vramData[13'd2775] = 8'd135;
vramData[13'd2776] = 8'd253;
vramData[13'd2777] = 8'd247;
vramData[13'd2778] = 8'd212;
vramData[13'd2779] = 8'd135;
vramData[13'd2780] = 8'd30;
vramData[13'd2781] = 8'd135;
vramData[13'd2782] = 8'd107;
vramData[13'd2783] = 8'd135;
vramData[13'd2784] = 8'd252;
vramData[13'd2785] = 8'd135;
vramData[13'd2786] = 8'd16;
vramData[13'd2787] = 8'd135;
vramData[13'd2788] = 8'd115;
vramData[13'd2789] = 8'd135;
vramData[13'd2790] = 8'd26;
vramData[13'd2791] = 8'd135;
vramData[13'd2792] = 8'd16;
vramData[13'd2793] = 8'd135;
vramData[13'd2794] = 8'd34;
vramData[13'd2795] = 8'd135;
vramData[13'd2796] = 8'd50;
vramData[13'd2797] = 8'd135;
vramData[13'd2798] = 8'd228;
vramData[13'd2799] = 8'd135;
vramData[13'd2800] = 8'd118;
vramData[13'd2801] = 8'd135;
vramData[13'd2802] = 8'd162;
vramData[13'd2803] = 8'd135;
vramData[13'd2804] = 8'd200;
vramData[13'd2805] = 8'd135;
vramData[13'd2806] = 8'd208;
vramData[13'd2807] = 8'd135;
vramData[13'd2808] = 8'd220;
vramData[13'd2809] = 8'd120;
vramData[13'd2810] = 8'd223;
vramData[13'd2811] = 8'd135;
vramData[13'd2812] = 8'd223;
vramData[13'd2813] = 8'd135;
vramData[13'd2814] = 8'd17;
vramData[13'd2815] = 8'd120;
vramData[13'd2816] = 8'd223;
vramData[13'd2817] = 8'd135;
vramData[13'd2818] = 8'd202;
vramData[13'd2819] = 8'd135;
vramData[13'd2820] = 8'd83;
vramData[13'd2821] = 8'd135;
vramData[13'd2822] = 8'd17;
vramData[13'd2823] = 8'd135;
vramData[13'd2824] = 8'd135;
vramData[13'd2825] = 8'd135;
vramData[13'd2826] = 8'd228;
vramData[13'd2827] = 8'd135;
vramData[13'd2828] = 8'd101;
vramData[13'd2829] = 8'd135;
vramData[13'd2830] = 8'd149;
vramData[13'd2831] = 8'd135;
vramData[13'd2832] = 8'd52;
vramData[13'd2833] = 8'd135;
vramData[13'd2834] = 8'd9;
vramData[13'd2835] = 8'd135;
vramData[13'd2836] = 8'd16;
vramData[13'd2837] = 8'd135;
vramData[13'd2838] = 8'd209;
vramData[13'd2839] = 8'd135;
vramData[13'd2840] = 8'd70;
vramData[13'd2841] = 8'd135;
vramData[13'd2842] = 8'd209;
vramData[13'd2843] = 8'd135;
vramData[13'd2844] = 8'd83;
vramData[13'd2845] = 8'd135;
vramData[13'd2846] = 8'd95;
vramData[13'd2847] = 8'd135;
vramData[13'd2848] = 8'd37;
vramData[13'd2849] = 8'd135;
vramData[13'd2850] = 8'd31;
vramData[13'd2851] = 8'd135;
vramData[13'd2852] = 8'd240;
vramData[13'd2853] = 8'd135;
vramData[13'd2854] = 8'd76;
vramData[13'd2855] = 8'd87;
vramData[13'd2856] = 8'd95;
vramData[13'd2857] = 8'd135;
vramData[13'd2858] = 8'd240;
vramData[13'd2859] = 8'd55;
vramData[13'd2860] = 8'd28;
vramData[13'd2861] = 8'd55;
vramData[13'd2862] = 8'd212;
vramData[13'd2863] = 8'd247;
vramData[13'd2864] = 8'd135;
vramData[13'd2865] = 8'd247;
vramData[13'd2866] = 8'd18;
vramData[13'd2867] = 8'd247;
vramData[13'd2868] = 8'd16;
vramData[13'd2869] = 8'd120;
vramData[13'd2870] = 8'd122;
vramData[13'd2871] = 8'd152;
vramData[13'd2872] = 8'd198;
vramData[13'd2873] = 8'd24;
vramData[13'd2874] = 8'd209;
vramData[13'd2875] = 8'd24;
vramData[13'd2876] = 8'd210;
vramData[13'd2877] = 8'd24;
vramData[13'd2878] = 8'd210;
vramData[13'd2879] = 8'd16;
vramData[13'd2880] = 8'd202;
vramData[13'd2881] = 8'd147;
vramData[13'd2882] = 8'd202;
vramData[13'd2883] = 8'd147;
vramData[13'd2884] = 8'd210;
vramData[13'd2885] = 8'd147;
vramData[13'd2886] = 8'd202;
vramData[13'd2887] = 8'd147;
vramData[13'd2888] = 8'd83;
vramData[13'd2889] = 8'd147;
vramData[13'd2890] = 8'd210;
vramData[13'd2891] = 8'd147;
vramData[13'd2892] = 8'd70;
vramData[13'd2893] = 8'd55;
vramData[13'd2894] = 8'd145;
vramData[13'd2895] = 8'd247;
vramData[13'd2896] = 8'd145;
vramData[13'd2897] = 8'd247;
vramData[13'd2898] = 8'd16;
vramData[13'd2899] = 8'd247;
vramData[13'd2900] = 8'd197;
vramData[13'd2901] = 8'd135;
vramData[13'd2902] = 8'd253;
vramData[13'd2903] = 8'd120;
vramData[13'd2904] = 8'd200;
vramData[13'd2905] = 8'd152;
vramData[13'd2906] = 8'd202;
vramData[13'd2907] = 8'd120;
vramData[13'd2908] = 8'd214;
vramData[13'd2909] = 8'd135;
vramData[13'd2910] = 8'd135;
vramData[13'd2911] = 8'd135;
vramData[13'd2912] = 8'd209;
vramData[13'd2913] = 8'd135;
vramData[13'd2914] = 8'd210;
vramData[13'd2915] = 8'd135;
vramData[13'd2916] = 8'd135;
vramData[13'd2917] = 8'd135;
vramData[13'd2918] = 8'd51;
vramData[13'd2919] = 8'd87;
vramData[13'd2920] = 8'd96;
vramData[13'd2921] = 8'd247;
vramData[13'd2922] = 8'd208;
vramData[13'd2923] = 8'd247;
vramData[13'd2924] = 8'd9;
vramData[13'd2925] = 8'd247;
vramData[13'd2926] = 8'd9;
vramData[13'd2927] = 8'd247;
vramData[13'd2928] = 8'd46;
vramData[13'd2929] = 8'd135;
vramData[13'd2930] = 8'd191;
vramData[13'd2931] = 8'd135;
vramData[13'd2932] = 8'd59;
vramData[13'd2933] = 8'd247;
vramData[13'd2934] = 8'd95;
vramData[13'd2935] = 8'd135;
vramData[13'd2936] = 8'd126;
vramData[13'd2937] = 8'd135;
vramData[13'd2938] = 8'd250;
vramData[13'd2939] = 8'd247;
vramData[13'd2940] = 8'd164;
vramData[13'd2941] = 8'd135;
vramData[13'd2942] = 8'd200;
vramData[13'd2943] = 8'd135;
vramData[13'd2944] = 8'd30;
vramData[13'd2945] = 8'd135;
vramData[13'd2946] = 8'd122;
vramData[13'd2947] = 8'd135;
vramData[13'd2948] = 8'd92;
vramData[13'd2949] = 8'd135;
vramData[13'd2950] = 8'd89;
vramData[13'd2951] = 8'd135;
vramData[13'd2952] = 8'd253;
vramData[13'd2953] = 8'd135;
vramData[13'd2954] = 8'd210;
vramData[13'd2955] = 8'd135;
vramData[13'd2956] = 8'd17;
vramData[13'd2957] = 8'd120;
vramData[13'd2958] = 8'd88;
vramData[13'd2959] = 8'd135;
vramData[13'd2960] = 8'd210;
vramData[13'd2961] = 8'd135;
vramData[13'd2962] = 8'd171;
vramData[13'd2963] = 8'd135;
vramData[13'd2964] = 8'd210;
vramData[13'd2965] = 8'd135;
vramData[13'd2966] = 8'd97;
vramData[13'd2967] = 8'd135;
vramData[13'd2968] = 8'd83;
vramData[13'd2969] = 8'd120;
vramData[13'd2970] = 8'd83;
vramData[13'd2971] = 8'd120;
vramData[13'd2972] = 8'd228;
vramData[13'd2973] = 8'd120;
vramData[13'd2974] = 8'd208;
vramData[13'd2975] = 8'd120;
vramData[13'd2976] = 8'd200;
vramData[13'd2977] = 8'd120;
vramData[13'd2978] = 8'd80;
vramData[13'd2979] = 8'd120;
vramData[13'd2980] = 8'd228;
vramData[13'd2981] = 8'd120;
vramData[13'd2982] = 8'd248;
vramData[13'd2983] = 8'd120;
vramData[13'd2984] = 8'd226;
vramData[13'd2985] = 8'd120;
vramData[13'd2986] = 8'd164;
vramData[13'd2987] = 8'd120;
vramData[13'd2988] = 8'd171;
vramData[13'd2989] = 8'd120;
vramData[13'd2990] = 8'd198;
vramData[13'd2991] = 8'd120;
vramData[13'd2992] = 8'd31;
vramData[13'd2993] = 8'd120;
vramData[13'd2994] = 8'd31;
vramData[13'd2995] = 8'd120;
vramData[13'd2996] = 8'd240;
vramData[13'd2997] = 8'd135;
vramData[13'd2998] = 8'd210;
vramData[13'd2999] = 8'd135;
vramData[13'd3000] = 8'd16;
vramData[13'd3001] = 8'd135;
vramData[13'd3002] = 8'd30;
vramData[13'd3003] = 8'd135;
vramData[13'd3004] = 8'd239;
vramData[13'd3005] = 8'd135;
vramData[13'd3006] = 8'd102;
vramData[13'd3007] = 8'd135;
vramData[13'd3008] = 8'd95;
vramData[13'd3009] = 8'd135;
vramData[13'd3010] = 8'd42;
vramData[13'd3011] = 8'd135;
vramData[13'd3012] = 8'd76;
vramData[13'd3013] = 8'd135;
vramData[13'd3014] = 8'd247;
vramData[13'd3015] = 8'd135;
vramData[13'd3016] = 8'd31;
vramData[13'd3017] = 8'd135;
vramData[13'd3018] = 8'd126;
vramData[13'd3019] = 8'd55;
vramData[13'd3020] = 8'd31;
vramData[13'd3021] = 8'd135;
vramData[13'd3022] = 8'd95;
vramData[13'd3023] = 8'd55;
vramData[13'd3024] = 8'd37;
vramData[13'd3025] = 8'd247;
vramData[13'd3026] = 8'd16;
vramData[13'd3027] = 8'd247;
vramData[13'd3028] = 8'd16;
vramData[13'd3029] = 8'd120;
vramData[13'd3030] = 8'd210;
vramData[13'd3031] = 8'd56;
vramData[13'd3032] = 8'd210;
vramData[13'd3033] = 8'd56;
vramData[13'd3034] = 8'd202;
vramData[13'd3035] = 8'd24;
vramData[13'd3036] = 8'd148;
vramData[13'd3037] = 8'd129;
vramData[13'd3038] = 8'd164;
vramData[13'd3039] = 8'd129;
vramData[13'd3040] = 8'd16;
vramData[13'd3041] = 8'd19;
vramData[13'd3042] = 8'd148;
vramData[13'd3043] = 8'd147;
vramData[13'd3044] = 8'd83;
vramData[13'd3045] = 8'd147;
vramData[13'd3046] = 8'd202;
vramData[13'd3047] = 8'd147;
vramData[13'd3048] = 8'd209;
vramData[13'd3049] = 8'd147;
vramData[13'd3050] = 8'd202;
vramData[13'd3051] = 8'd147;
vramData[13'd3052] = 8'd135;
vramData[13'd3053] = 8'd55;
vramData[13'd3054] = 8'd214;
vramData[13'd3055] = 8'd55;
vramData[13'd3056] = 8'd95;
vramData[13'd3057] = 8'd135;
vramData[13'd3058] = 8'd210;
vramData[13'd3059] = 8'd135;
vramData[13'd3060] = 8'd155;
vramData[13'd3061] = 8'd135;
vramData[13'd3062] = 8'd16;
vramData[13'd3063] = 8'd120;
vramData[13'd3064] = 8'd108;
vramData[13'd3065] = 8'd8;
vramData[13'd3066] = 8'd96;
vramData[13'd3067] = 8'd8;
vramData[13'd3068] = 8'd214;
vramData[13'd3069] = 8'd8;
vramData[13'd3070] = 8'd94;
vramData[13'd3071] = 8'd120;
vramData[13'd3072] = 8'd252;
vramData[13'd3073] = 8'd152;
vramData[13'd3074] = 8'd252;
vramData[13'd3075] = 8'd152;
vramData[13'd3076] = 8'd200;
vramData[13'd3077] = 8'd120;
vramData[13'd3078] = 8'd16;
vramData[13'd3079] = 8'd135;
vramData[13'd3080] = 8'd110;
vramData[13'd3081] = 8'd247;
vramData[13'd3082] = 8'd219;
vramData[13'd3083] = 8'd123;
vramData[13'd3084] = 8'd96;
vramData[13'd3085] = 8'd247;
vramData[13'd3086] = 8'd196;
vramData[13'd3087] = 8'd247;
vramData[13'd3088] = 8'd30;
vramData[13'd3089] = 8'd87;
vramData[13'd3090] = 8'd93;
vramData[13'd3091] = 8'd135;
vramData[13'd3092] = 8'd116;
vramData[13'd3093] = 8'd119;
vramData[13'd3094] = 8'd17;
vramData[13'd3095] = 8'd247;
vramData[13'd3096] = 8'd251;
vramData[13'd3097] = 8'd247;
vramData[13'd3098] = 8'd16;
vramData[13'd3099] = 8'd247;
vramData[13'd3100] = 8'd251;
vramData[13'd3101] = 8'd135;
vramData[13'd3102] = 8'd210;
vramData[13'd3103] = 8'd135;
vramData[13'd3104] = 8'd37;
vramData[13'd3105] = 8'd135;
vramData[13'd3106] = 8'd244;
vramData[13'd3107] = 8'd135;
vramData[13'd3108] = 8'd101;
vramData[13'd3109] = 8'd135;
vramData[13'd3110] = 8'd30;
vramData[13'd3111] = 8'd135;
vramData[13'd3112] = 8'd97;
vramData[13'd3113] = 8'd135;
vramData[13'd3114] = 8'd148;
vramData[13'd3115] = 8'd120;
vramData[13'd3116] = 8'd30;
vramData[13'd3117] = 8'd120;
vramData[13'd3118] = 8'd83;
vramData[13'd3119] = 8'd120;
vramData[13'd3120] = 8'd135;
vramData[13'd3121] = 8'd120;
vramData[13'd3122] = 8'd164;
vramData[13'd3123] = 8'd120;
vramData[13'd3124] = 8'd210;
vramData[13'd3125] = 8'd120;
vramData[13'd3126] = 8'd155;
vramData[13'd3127] = 8'd120;
vramData[13'd3128] = 8'd202;
vramData[13'd3129] = 8'd135;
vramData[13'd3130] = 8'd30;
vramData[13'd3131] = 8'd120;
vramData[13'd3132] = 8'd70;
vramData[13'd3133] = 8'd120;
vramData[13'd3134] = 8'd135;
vramData[13'd3135] = 8'd120;
vramData[13'd3136] = 8'd135;
vramData[13'd3137] = 8'd120;
vramData[13'd3138] = 8'd30;
vramData[13'd3139] = 8'd120;
vramData[13'd3140] = 8'd18;
vramData[13'd3141] = 8'd152;
vramData[13'd3142] = 8'd214;
vramData[13'd3143] = 8'd120;
vramData[13'd3144] = 8'd240;
vramData[13'd3145] = 8'd120;
vramData[13'd3146] = 8'd210;
vramData[13'd3147] = 8'd120;
vramData[13'd3148] = 8'd17;
vramData[13'd3149] = 8'd120;
vramData[13'd3150] = 8'd101;
vramData[13'd3151] = 8'd120;
vramData[13'd3152] = 8'd214;
vramData[13'd3153] = 8'd120;
vramData[13'd3154] = 8'd80;
vramData[13'd3155] = 8'd135;
vramData[13'd3156] = 8'd115;
vramData[13'd3157] = 8'd135;
vramData[13'd3158] = 8'd70;
vramData[13'd3159] = 8'd135;
vramData[13'd3160] = 8'd31;
vramData[13'd3161] = 8'd135;
vramData[13'd3162] = 8'd31;
vramData[13'd3163] = 8'd135;
vramData[13'd3164] = 8'd94;
vramData[13'd3165] = 8'd135;
vramData[13'd3166] = 8'd248;
vramData[13'd3167] = 8'd135;
vramData[13'd3168] = 8'd92;
vramData[13'd3169] = 8'd135;
vramData[13'd3170] = 8'd83;
vramData[13'd3171] = 8'd135;
vramData[13'd3172] = 8'd200;
vramData[13'd3173] = 8'd135;
vramData[13'd3174] = 8'd80;
vramData[13'd3175] = 8'd87;
vramData[13'd3176] = 8'd184;
vramData[13'd3177] = 8'd135;
vramData[13'd3178] = 8'd28;
vramData[13'd3179] = 8'd87;
vramData[13'd3180] = 8'd29;
vramData[13'd3181] = 8'd247;
vramData[13'd3182] = 8'd95;
vramData[13'd3183] = 8'd247;
vramData[13'd3184] = 8'd200;
vramData[13'd3185] = 8'd247;
vramData[13'd3186] = 8'd16;
vramData[13'd3187] = 8'd247;
vramData[13'd3188] = 8'd198;
vramData[13'd3189] = 8'd55;
vramData[13'd3190] = 8'd16;
vramData[13'd3191] = 8'd115;
vramData[13'd3192] = 8'd210;
vramData[13'd3193] = 8'd115;
vramData[13'd3194] = 8'd202;
vramData[13'd3195] = 8'd147;
vramData[13'd3196] = 8'd202;
vramData[13'd3197] = 8'd19;
vramData[13'd3198] = 8'd210;
vramData[13'd3199] = 8'd49;
vramData[13'd3200] = 8'd202;
vramData[13'd3201] = 8'd56;
vramData[13'd3202] = 8'd210;
vramData[13'd3203] = 8'd131;
vramData[13'd3204] = 8'd202;
vramData[13'd3205] = 8'd147;
vramData[13'd3206] = 8'd202;
vramData[13'd3207] = 8'd147;
vramData[13'd3208] = 8'd202;
vramData[13'd3209] = 8'd147;
vramData[13'd3210] = 8'd80;
vramData[13'd3211] = 8'd147;
vramData[13'd3212] = 8'd80;
vramData[13'd3213] = 8'd147;
vramData[13'd3214] = 8'd16;
vramData[13'd3215] = 8'd55;
vramData[13'd3216] = 8'd80;
vramData[13'd3217] = 8'd135;
vramData[13'd3218] = 8'd226;
vramData[13'd3219] = 8'd135;
vramData[13'd3220] = 8'd228;
vramData[13'd3221] = 8'd135;
vramData[13'd3222] = 8'd0;
vramData[13'd3223] = 8'd199;
vramData[13'd3224] = 8'd16;
vramData[13'd3225] = 8'd120;
vramData[13'd3226] = 8'd209;
vramData[13'd3227] = 8'd8;
vramData[13'd3228] = 8'd16;
vramData[13'd3229] = 8'd8;
vramData[13'd3230] = 8'd81;
vramData[13'd3231] = 8'd136;
vramData[13'd3232] = 8'd95;
vramData[13'd3233] = 8'd8;
vramData[13'd3234] = 8'd183;
vramData[13'd3235] = 8'd8;
vramData[13'd3236] = 8'd95;
vramData[13'd3237] = 8'd8;
vramData[13'd3238] = 8'd94;
vramData[13'd3239] = 8'd120;
vramData[13'd3240] = 8'd223;
vramData[13'd3241] = 8'd120;
vramData[13'd3242] = 8'd223;
vramData[13'd3243] = 8'd120;
vramData[13'd3244] = 8'd183;
vramData[13'd3245] = 8'd135;
vramData[13'd3246] = 8'd210;
vramData[13'd3247] = 8'd135;
vramData[13'd3248] = 8'd230;
vramData[13'd3249] = 8'd135;
vramData[13'd3250] = 8'd31;
vramData[13'd3251] = 8'd247;
vramData[13'd3252] = 8'd208;
vramData[13'd3253] = 8'd247;
vramData[13'd3254] = 8'd248;
vramData[13'd3255] = 8'd247;
vramData[13'd3256] = 8'd200;
vramData[13'd3257] = 8'd247;
vramData[13'd3258] = 8'd155;
vramData[13'd3259] = 8'd247;
vramData[13'd3260] = 8'd28;
vramData[13'd3261] = 8'd247;
vramData[13'd3262] = 8'd155;
vramData[13'd3263] = 8'd135;
vramData[13'd3264] = 8'd149;
vramData[13'd3265] = 8'd135;
vramData[13'd3266] = 8'd240;
vramData[13'd3267] = 8'd135;
vramData[13'd3268] = 8'd31;
vramData[13'd3269] = 8'd135;
vramData[13'd3270] = 8'd101;
vramData[13'd3271] = 8'd120;
vramData[13'd3272] = 8'd135;
vramData[13'd3273] = 8'd135;
vramData[13'd3274] = 8'd90;
vramData[13'd3275] = 8'd135;
vramData[13'd3276] = 8'd156;
vramData[13'd3277] = 8'd135;
vramData[13'd3278] = 8'd155;
vramData[13'd3279] = 8'd120;
vramData[13'd3280] = 8'd37;
vramData[13'd3281] = 8'd120;
vramData[13'd3282] = 8'd156;
vramData[13'd3283] = 8'd120;
vramData[13'd3284] = 8'd202;
vramData[13'd3285] = 8'd120;
vramData[13'd3286] = 8'd83;
vramData[13'd3287] = 8'd120;
vramData[13'd3288] = 8'd17;
vramData[13'd3289] = 8'd120;
vramData[13'd3290] = 8'd145;
vramData[13'd3291] = 8'd120;
vramData[13'd3292] = 8'd30;
vramData[13'd3293] = 8'd120;
vramData[13'd3294] = 8'd101;
vramData[13'd3295] = 8'd120;
vramData[13'd3296] = 8'd202;
vramData[13'd3297] = 8'd120;
vramData[13'd3298] = 8'd30;
vramData[13'd3299] = 8'd120;
vramData[13'd3300] = 8'd83;
vramData[13'd3301] = 8'd120;
vramData[13'd3302] = 8'd83;
vramData[13'd3303] = 8'd120;
vramData[13'd3304] = 8'd30;
vramData[13'd3305] = 8'd120;
vramData[13'd3306] = 8'd80;
vramData[13'd3307] = 8'd135;
vramData[13'd3308] = 8'd80;
vramData[13'd3309] = 8'd120;
vramData[13'd3310] = 8'd164;
vramData[13'd3311] = 8'd135;
vramData[13'd3312] = 8'd31;
vramData[13'd3313] = 8'd135;
vramData[13'd3314] = 8'd16;
vramData[13'd3315] = 8'd135;
vramData[13'd3316] = 8'd200;
vramData[13'd3317] = 8'd135;
vramData[13'd3318] = 8'd17;
vramData[13'd3319] = 8'd135;
vramData[13'd3320] = 8'd248;
vramData[13'd3321] = 8'd135;
vramData[13'd3322] = 8'd253;
vramData[13'd3323] = 8'd103;
vramData[13'd3324] = 8'd150;
vramData[13'd3325] = 8'd119;
vramData[13'd3326] = 8'd251;
vramData[13'd3327] = 8'd55;
vramData[13'd3328] = 8'd83;
vramData[13'd3329] = 8'd135;
vramData[13'd3330] = 8'd249;
vramData[13'd3331] = 8'd135;
vramData[13'd3332] = 8'd31;
vramData[13'd3333] = 8'd135;
vramData[13'd3334] = 8'd31;
vramData[13'd3335] = 8'd135;
vramData[13'd3336] = 8'd191;
vramData[13'd3337] = 8'd135;
vramData[13'd3338] = 8'd170;
vramData[13'd3339] = 8'd247;
vramData[13'd3340] = 8'd95;
vramData[13'd3341] = 8'd247;
vramData[13'd3342] = 8'd198;
vramData[13'd3343] = 8'd247;
vramData[13'd3344] = 8'd202;
vramData[13'd3345] = 8'd247;
vramData[13'd3346] = 8'd16;
vramData[13'd3347] = 8'd247;
vramData[13'd3348] = 8'd80;
vramData[13'd3349] = 8'd115;
vramData[13'd3350] = 8'd31;
vramData[13'd3351] = 8'd147;
vramData[13'd3352] = 8'd16;
vramData[13'd3353] = 8'd147;
vramData[13'd3354] = 8'd210;
vramData[13'd3355] = 8'd19;
vramData[13'd3356] = 8'd210;
vramData[13'd3357] = 8'd131;
vramData[13'd3358] = 8'd210;
vramData[13'd3359] = 8'd131;
vramData[13'd3360] = 8'd202;
vramData[13'd3361] = 8'd24;
vramData[13'd3362] = 8'd202;
vramData[13'd3363] = 8'd56;
vramData[13'd3364] = 8'd145;
vramData[13'd3365] = 8'd56;
vramData[13'd3366] = 8'd16;
vramData[13'd3367] = 8'd56;
vramData[13'd3368] = 8'd202;
vramData[13'd3369] = 8'd24;
vramData[13'd3370] = 8'd37;
vramData[13'd3371] = 8'd8;
vramData[13'd3372] = 8'd16;
vramData[13'd3373] = 8'd8;
vramData[13'd3374] = 8'd198;
vramData[13'd3375] = 8'd152;
vramData[13'd3376] = 8'd37;
vramData[13'd3377] = 8'd135;
vramData[13'd3378] = 8'd16;
vramData[13'd3379] = 8'd135;
vramData[13'd3380] = 8'd16;
vramData[13'd3381] = 8'd135;
vramData[13'd3382] = 8'd166;
vramData[13'd3383] = 8'd87;
vramData[13'd3384] = 8'd221;
vramData[13'd3385] = 8'd120;
vramData[13'd3386] = 8'd202;
vramData[13'd3387] = 8'd8;
vramData[13'd3388] = 8'd16;
vramData[13'd3389] = 8'd8;
vramData[13'd3390] = 8'd52;
vramData[13'd3391] = 8'd200;
vramData[13'd3392] = 8'd168;
vramData[13'd3393] = 8'd120;
vramData[13'd3394] = 8'd198;
vramData[13'd3395] = 8'd8;
vramData[13'd3396] = 8'd80;
vramData[13'd3397] = 8'd8;
vramData[13'd3398] = 8'd95;
vramData[13'd3399] = 8'd120;
vramData[13'd3400] = 8'd214;
vramData[13'd3401] = 8'd120;
vramData[13'd3402] = 8'd214;
vramData[13'd3403] = 8'd120;
vramData[13'd3404] = 8'd223;
vramData[13'd3405] = 8'd135;
vramData[13'd3406] = 8'd252;
vramData[13'd3407] = 8'd135;
vramData[13'd3408] = 8'd60;
vramData[13'd3409] = 8'd247;
vramData[13'd3410] = 8'd243;
vramData[13'd3411] = 8'd247;
vramData[13'd3412] = 8'd18;
vramData[13'd3413] = 8'd247;
vramData[13'd3414] = 8'd240;
vramData[13'd3415] = 8'd247;
vramData[13'd3416] = 8'd212;
vramData[13'd3417] = 8'd247;
vramData[13'd3418] = 8'd166;
vramData[13'd3419] = 8'd135;
vramData[13'd3420] = 8'd210;
vramData[13'd3421] = 8'd135;
vramData[13'd3422] = 8'd135;
vramData[13'd3423] = 8'd135;
vramData[13'd3424] = 8'd67;
vramData[13'd3425] = 8'd135;
vramData[13'd3426] = 8'd122;
vramData[13'd3427] = 8'd135;
vramData[13'd3428] = 8'd209;
vramData[13'd3429] = 8'd135;
vramData[13'd3430] = 8'd83;
vramData[13'd3431] = 8'd135;
vramData[13'd3432] = 8'd228;
vramData[13'd3433] = 8'd120;
vramData[13'd3434] = 8'd31;
vramData[13'd3435] = 8'd135;
vramData[13'd3436] = 8'd202;
vramData[13'd3437] = 8'd135;
vramData[13'd3438] = 8'd31;
vramData[13'd3439] = 8'd135;
vramData[13'd3440] = 8'd80;
vramData[13'd3441] = 8'd120;
vramData[13'd3442] = 8'd208;
vramData[13'd3443] = 8'd120;
vramData[13'd3444] = 8'd240;
vramData[13'd3445] = 8'd120;
vramData[13'd3446] = 8'd205;
vramData[13'd3447] = 8'd120;
vramData[13'd3448] = 8'd239;
vramData[13'd3449] = 8'd120;
vramData[13'd3450] = 8'd31;
vramData[13'd3451] = 8'd120;
vramData[13'd3452] = 8'd30;
vramData[13'd3453] = 8'd120;
vramData[13'd3454] = 8'd31;
vramData[13'd3455] = 8'd120;
vramData[13'd3456] = 8'd31;
vramData[13'd3457] = 8'd120;
vramData[13'd3458] = 8'd239;
vramData[13'd3459] = 8'd120;
vramData[13'd3460] = 8'd83;
vramData[13'd3461] = 8'd120;
vramData[13'd3462] = 8'd37;
vramData[13'd3463] = 8'd120;
vramData[13'd3464] = 8'd240;
vramData[13'd3465] = 8'd135;
vramData[13'd3466] = 8'd31;
vramData[13'd3467] = 8'd135;
vramData[13'd3468] = 8'd30;
vramData[13'd3469] = 8'd135;
vramData[13'd3470] = 8'd145;
vramData[13'd3471] = 8'd135;
vramData[13'd3472] = 8'd156;
vramData[13'd3473] = 8'd135;
vramData[13'd3474] = 8'd90;
vramData[13'd3475] = 8'd135;
vramData[13'd3476] = 8'd95;
vramData[13'd3477] = 8'd135;
vramData[13'd3478] = 8'd115;
vramData[13'd3479] = 8'd135;
vramData[13'd3480] = 8'd67;
vramData[13'd3481] = 8'd135;
vramData[13'd3482] = 8'd228;
vramData[13'd3483] = 8'd135;
vramData[13'd3484] = 8'd95;
vramData[13'd3485] = 8'd135;
vramData[13'd3486] = 8'd31;
vramData[13'd3487] = 8'd135;
vramData[13'd3488] = 8'd29;
vramData[13'd3489] = 8'd135;
vramData[13'd3490] = 8'd135;
vramData[13'd3491] = 8'd135;
vramData[13'd3492] = 8'd190;
vramData[13'd3493] = 8'd135;
vramData[13'd3494] = 8'd211;
vramData[13'd3495] = 8'd135;
vramData[13'd3496] = 8'd248;
vramData[13'd3497] = 8'd135;
vramData[13'd3498] = 8'd170;
vramData[13'd3499] = 8'd247;
vramData[13'd3500] = 8'd50;
vramData[13'd3501] = 8'd247;
vramData[13'd3502] = 8'd30;
vramData[13'd3503] = 8'd247;
vramData[13'd3504] = 8'd210;
vramData[13'd3505] = 8'd247;
vramData[13'd3506] = 8'd16;
vramData[13'd3507] = 8'd247;
vramData[13'd3508] = 8'd16;
vramData[13'd3509] = 8'd115;
vramData[13'd3510] = 8'd210;
vramData[13'd3511] = 8'd131;
vramData[13'd3512] = 8'd210;
vramData[13'd3513] = 8'd131;
vramData[13'd3514] = 8'd202;
vramData[13'd3515] = 8'd56;
vramData[13'd3516] = 8'd209;
vramData[13'd3517] = 8'd56;
vramData[13'd3518] = 8'd209;
vramData[13'd3519] = 8'd56;
vramData[13'd3520] = 8'd210;
vramData[13'd3521] = 8'd24;
vramData[13'd3522] = 8'd210;
vramData[13'd3523] = 8'd24;
vramData[13'd3524] = 8'd202;
vramData[13'd3525] = 8'd56;
vramData[13'd3526] = 8'd148;
vramData[13'd3527] = 8'd56;
vramData[13'd3528] = 8'd16;
vramData[13'd3529] = 8'd56;
vramData[13'd3530] = 8'd127;
vramData[13'd3531] = 8'd120;
vramData[13'd3532] = 8'd30;
vramData[13'd3533] = 8'd120;
vramData[13'd3534] = 8'd31;
vramData[13'd3535] = 8'd120;
vramData[13'd3536] = 8'd200;
vramData[13'd3537] = 8'd120;
vramData[13'd3538] = 8'd210;
vramData[13'd3539] = 8'd135;
vramData[13'd3540] = 8'd210;
vramData[13'd3541] = 8'd135;
vramData[13'd3542] = 8'd16;
vramData[13'd3543] = 8'd135;
vramData[13'd3544] = 8'd212;
vramData[13'd3545] = 8'd55;
vramData[13'd3546] = 8'd16;
vramData[13'd3547] = 8'd120;
vramData[13'd3548] = 8'd83;
vramData[13'd3549] = 8'd8;
vramData[13'd3550] = 8'd80;
vramData[13'd3551] = 8'd8;
vramData[13'd3552] = 8'd16;
vramData[13'd3553] = 8'd8;
vramData[13'd3554] = 8'd172;
vramData[13'd3555] = 8'd120;
vramData[13'd3556] = 8'd164;
vramData[13'd3557] = 8'd135;
vramData[13'd3558] = 8'd94;
vramData[13'd3559] = 8'd135;
vramData[13'd3560] = 8'd141;
vramData[13'd3561] = 8'd135;
vramData[13'd3562] = 8'd145;
vramData[13'd3563] = 8'd247;
vramData[13'd3564] = 8'd139;
vramData[13'd3565] = 8'd247;
vramData[13'd3566] = 8'd211;
vramData[13'd3567] = 8'd247;
vramData[13'd3568] = 8'd45;
vramData[13'd3569] = 8'd135;
vramData[13'd3570] = 8'd46;
vramData[13'd3571] = 8'd135;
vramData[13'd3572] = 8'd192;
vramData[13'd3573] = 8'd247;
vramData[13'd3574] = 8'd92;
vramData[13'd3575] = 8'd135;
vramData[13'd3576] = 8'd127;
vramData[13'd3577] = 8'd135;
vramData[13'd3578] = 8'd218;
vramData[13'd3579] = 8'd135;
vramData[13'd3580] = 8'd200;
vramData[13'd3581] = 8'd135;
vramData[13'd3582] = 8'd240;
vramData[13'd3583] = 8'd135;
vramData[13'd3584] = 8'd9;
vramData[13'd3585] = 8'd135;
vramData[13'd3586] = 8'd230;
vramData[13'd3587] = 8'd135;
vramData[13'd3588] = 8'd164;
vramData[13'd3589] = 8'd135;
vramData[13'd3590] = 8'd240;
vramData[13'd3591] = 8'd120;
vramData[13'd3592] = 8'd83;
vramData[13'd3593] = 8'd120;
vramData[13'd3594] = 8'd90;
vramData[13'd3595] = 8'd120;
vramData[13'd3596] = 8'd42;
vramData[13'd3597] = 8'd120;
vramData[13'd3598] = 8'd16;
vramData[13'd3599] = 8'd135;
vramData[13'd3600] = 8'd240;
vramData[13'd3601] = 8'd120;
vramData[13'd3602] = 8'd30;
vramData[13'd3603] = 8'd135;
vramData[13'd3604] = 8'd115;
vramData[13'd3605] = 8'd120;
vramData[13'd3606] = 8'd122;
vramData[13'd3607] = 8'd120;
vramData[13'd3608] = 8'd240;
vramData[13'd3609] = 8'd120;
vramData[13'd3610] = 8'd31;
vramData[13'd3611] = 8'd120;
vramData[13'd3612] = 8'd30;
vramData[13'd3613] = 8'd120;
vramData[13'd3614] = 8'd83;
vramData[13'd3615] = 8'd120;
vramData[13'd3616] = 8'd155;
vramData[13'd3617] = 8'd120;
vramData[13'd3618] = 8'd211;
vramData[13'd3619] = 8'd120;
vramData[13'd3620] = 8'd83;
vramData[13'd3621] = 8'd120;
vramData[13'd3622] = 8'd80;
vramData[13'd3623] = 8'd135;
vramData[13'd3624] = 8'd80;
vramData[13'd3625] = 8'd135;
vramData[13'd3626] = 8'd30;
vramData[13'd3627] = 8'd135;
vramData[13'd3628] = 8'd90;
vramData[13'd3629] = 8'd135;
vramData[13'd3630] = 8'd210;
vramData[13'd3631] = 8'd135;
vramData[13'd3632] = 8'd50;
vramData[13'd3633] = 8'd135;
vramData[13'd3634] = 8'd37;
vramData[13'd3635] = 8'd135;
vramData[13'd3636] = 8'd135;
vramData[13'd3637] = 8'd135;
vramData[13'd3638] = 8'd31;
vramData[13'd3639] = 8'd135;
vramData[13'd3640] = 8'd251;
vramData[13'd3641] = 8'd135;
vramData[13'd3642] = 8'd90;
vramData[13'd3643] = 8'd135;
vramData[13'd3644] = 8'd30;
vramData[13'd3645] = 8'd135;
vramData[13'd3646] = 8'd228;
vramData[13'd3647] = 8'd55;
vramData[13'd3648] = 8'd248;
vramData[13'd3649] = 8'd135;
vramData[13'd3650] = 8'd207;
vramData[13'd3651] = 8'd135;
vramData[13'd3652] = 8'd51;
vramData[13'd3653] = 8'd135;
vramData[13'd3654] = 8'd28;
vramData[13'd3655] = 8'd135;
vramData[13'd3656] = 8'd96;
vramData[13'd3657] = 8'd135;
vramData[13'd3658] = 8'd95;
vramData[13'd3659] = 8'd247;
vramData[13'd3660] = 8'd30;
vramData[13'd3661] = 8'd247;
vramData[13'd3662] = 8'd148;
vramData[13'd3663] = 8'd247;
vramData[13'd3664] = 8'd16;
vramData[13'd3665] = 8'd247;
vramData[13'd3666] = 8'd198;
vramData[13'd3667] = 8'd55;
vramData[13'd3668] = 8'd16;
vramData[13'd3669] = 8'd115;
vramData[13'd3670] = 8'd210;
vramData[13'd3671] = 8'd147;
vramData[13'd3672] = 8'd210;
vramData[13'd3673] = 8'd147;
vramData[13'd3674] = 8'd202;
vramData[13'd3675] = 8'd19;
vramData[13'd3676] = 8'd202;
vramData[13'd3677] = 8'd19;
vramData[13'd3678] = 8'd202;
vramData[13'd3679] = 8'd19;
vramData[13'd3680] = 8'd202;
vramData[13'd3681] = 8'd24;
vramData[13'd3682] = 8'd202;
vramData[13'd3683] = 8'd24;
vramData[13'd3684] = 8'd202;
vramData[13'd3685] = 8'd152;
vramData[13'd3686] = 8'd202;
vramData[13'd3687] = 8'd56;
vramData[13'd3688] = 8'd202;
vramData[13'd3689] = 8'd152;
vramData[13'd3690] = 8'd210;
vramData[13'd3691] = 8'd152;
vramData[13'd3692] = 8'd210;
vramData[13'd3693] = 8'd152;
vramData[13'd3694] = 8'd135;
vramData[13'd3695] = 8'd152;
vramData[13'd3696] = 8'd214;
vramData[13'd3697] = 8'd152;
vramData[13'd3698] = 8'd210;
vramData[13'd3699] = 8'd120;
vramData[13'd3700] = 8'd209;
vramData[13'd3701] = 8'd120;
vramData[13'd3702] = 8'd80;
vramData[13'd3703] = 8'd135;
vramData[13'd3704] = 8'd214;
vramData[13'd3705] = 8'd135;
vramData[13'd3706] = 8'd16;
vramData[13'd3707] = 8'd120;
vramData[13'd3708] = 8'd117;
vramData[13'd3709] = 8'd152;
vramData[13'd3710] = 8'd45;
vramData[13'd3711] = 8'd8;
vramData[13'd3712] = 8'd88;
vramData[13'd3713] = 8'd120;
vramData[13'd3714] = 8'd95;
vramData[13'd3715] = 8'd135;
vramData[13'd3716] = 8'd252;
vramData[13'd3717] = 8'd135;
vramData[13'd3718] = 8'd247;
vramData[13'd3719] = 8'd247;
vramData[13'd3720] = 8'd94;
vramData[13'd3721] = 8'd135;
vramData[13'd3722] = 8'd62;
vramData[13'd3723] = 8'd135;
vramData[13'd3724] = 8'd46;
vramData[13'd3725] = 8'd135;
vramData[13'd3726] = 8'd252;
vramData[13'd3727] = 8'd135;
vramData[13'd3728] = 8'd96;
vramData[13'd3729] = 8'd247;
vramData[13'd3730] = 8'd30;
vramData[13'd3731] = 8'd135;
vramData[13'd3732] = 8'd16;
vramData[13'd3733] = 8'd135;
vramData[13'd3734] = 8'd149;
vramData[13'd3735] = 8'd135;
vramData[13'd3736] = 8'd171;
vramData[13'd3737] = 8'd120;
vramData[13'd3738] = 8'd51;
vramData[13'd3739] = 8'd120;
vramData[13'd3740] = 8'd85;
vramData[13'd3741] = 8'd135;
vramData[13'd3742] = 8'd200;
vramData[13'd3743] = 8'd120;
vramData[13'd3744] = 8'd83;
vramData[13'd3745] = 8'd135;
vramData[13'd3746] = 8'd55;
vramData[13'd3747] = 8'd135;
vramData[13'd3748] = 8'd9;
vramData[13'd3749] = 8'd120;
vramData[13'd3750] = 8'd164;
vramData[13'd3751] = 8'd135;
vramData[13'd3752] = 8'd83;
vramData[13'd3753] = 8'd120;
vramData[13'd3754] = 8'd166;
vramData[13'd3755] = 8'd120;
vramData[13'd3756] = 8'd31;
vramData[13'd3757] = 8'd120;
vramData[13'd3758] = 8'd115;
vramData[13'd3759] = 8'd120;
vramData[13'd3760] = 8'd16;
vramData[13'd3761] = 8'd135;
vramData[13'd3762] = 8'd171;
vramData[13'd3763] = 8'd135;
vramData[13'd3764] = 8'd208;
vramData[13'd3765] = 8'd135;
vramData[13'd3766] = 8'd31;
vramData[13'd3767] = 8'd120;
vramData[13'd3768] = 8'd145;
vramData[13'd3769] = 8'd120;
vramData[13'd3770] = 8'd30;
vramData[13'd3771] = 8'd120;
vramData[13'd3772] = 8'd135;
vramData[13'd3773] = 8'd120;
vramData[13'd3774] = 8'd16;
vramData[13'd3775] = 8'd120;
vramData[13'd3776] = 8'd135;
vramData[13'd3777] = 8'd120;
vramData[13'd3778] = 8'd210;
vramData[13'd3779] = 8'd120;
vramData[13'd3780] = 8'd31;
vramData[13'd3781] = 8'd135;
vramData[13'd3782] = 8'd148;
vramData[13'd3783] = 8'd120;
vramData[13'd3784] = 8'd164;
vramData[13'd3785] = 8'd120;
vramData[13'd3786] = 8'd80;
vramData[13'd3787] = 8'd120;
vramData[13'd3788] = 8'd228;
vramData[13'd3789] = 8'd120;
vramData[13'd3790] = 8'd200;
vramData[13'd3791] = 8'd120;
vramData[13'd3792] = 8'd145;
vramData[13'd3793] = 8'd135;
vramData[13'd3794] = 8'd95;
vramData[13'd3795] = 8'd135;
vramData[13'd3796] = 8'd90;
vramData[13'd3797] = 8'd135;
vramData[13'd3798] = 8'd210;
vramData[13'd3799] = 8'd135;
vramData[13'd3800] = 8'd238;
vramData[13'd3801] = 8'd135;
vramData[13'd3802] = 8'd91;
vramData[13'd3803] = 8'd135;
vramData[13'd3804] = 8'd240;
vramData[13'd3805] = 8'd135;
vramData[13'd3806] = 8'd229;
vramData[13'd3807] = 8'd55;
vramData[13'd3808] = 8'd90;
vramData[13'd3809] = 8'd55;
vramData[13'd3810] = 8'd250;
vramData[13'd3811] = 8'd135;
vramData[13'd3812] = 8'd30;
vramData[13'd3813] = 8'd135;
vramData[13'd3814] = 8'd228;
vramData[13'd3815] = 8'd135;
vramData[13'd3816] = 8'd116;
vramData[13'd3817] = 8'd87;
vramData[13'd3818] = 8'd148;
vramData[13'd3819] = 8'd119;
vramData[13'd3820] = 8'd95;
vramData[13'd3821] = 8'd247;
vramData[13'd3822] = 8'd80;
vramData[13'd3823] = 8'd247;
vramData[13'd3824] = 8'd235;
vramData[13'd3825] = 8'd119;
vramData[13'd3826] = 8'd198;
vramData[13'd3827] = 8'd183;
vramData[13'd3828] = 8'd80;
vramData[13'd3829] = 8'd123;
vramData[13'd3830] = 8'd210;
vramData[13'd3831] = 8'd179;
vramData[13'd3832] = 8'd210;
vramData[13'd3833] = 8'd179;
vramData[13'd3834] = 8'd210;
vramData[13'd3835] = 8'd179;
vramData[13'd3836] = 8'd210;
vramData[13'd3837] = 8'd179;
vramData[13'd3838] = 8'd210;
vramData[13'd3839] = 8'd147;
vramData[13'd3840] = 8'd209;
vramData[13'd3841] = 8'd152;
vramData[13'd3842] = 8'd164;
vramData[13'd3843] = 8'd152;
vramData[13'd3844] = 8'd83;
vramData[13'd3845] = 8'd152;
vramData[13'd3846] = 8'd30;
vramData[13'd3847] = 8'd152;
vramData[13'd3848] = 8'd181;
vramData[13'd3849] = 8'd152;
vramData[13'd3850] = 8'd145;
vramData[13'd3851] = 8'd152;
vramData[13'd3852] = 8'd210;
vramData[13'd3853] = 8'd152;
vramData[13'd3854] = 8'd148;
vramData[13'd3855] = 8'd152;
vramData[13'd3856] = 8'd31;
vramData[13'd3857] = 8'd120;
vramData[13'd3858] = 8'd80;
vramData[13'd3859] = 8'd120;
vramData[13'd3860] = 8'd210;
vramData[13'd3861] = 8'd152;
vramData[13'd3862] = 8'd202;
vramData[13'd3863] = 8'd120;
vramData[13'd3864] = 8'd210;
vramData[13'd3865] = 8'd135;
vramData[13'd3866] = 8'd202;
vramData[13'd3867] = 8'd120;
vramData[13'd3868] = 8'd31;
vramData[13'd3869] = 8'd152;
vramData[13'd3870] = 8'd16;
vramData[13'd3871] = 8'd152;
vramData[13'd3872] = 8'd104;
vramData[13'd3873] = 8'd120;
vramData[13'd3874] = 8'd164;
vramData[13'd3875] = 8'd120;
vramData[13'd3876] = 8'd198;
vramData[13'd3877] = 8'd120;
vramData[13'd3878] = 8'd135;
vramData[13'd3879] = 8'd135;
vramData[13'd3880] = 8'd244;
vramData[13'd3881] = 8'd135;
vramData[13'd3882] = 8'd107;
vramData[13'd3883] = 8'd135;
vramData[13'd3884] = 8'd230;
vramData[13'd3885] = 8'd135;
vramData[13'd3886] = 8'd200;
vramData[13'd3887] = 8'd135;
vramData[13'd3888] = 8'd248;
vramData[13'd3889] = 8'd120;
vramData[13'd3890] = 8'd16;
vramData[13'd3891] = 8'd135;
vramData[13'd3892] = 8'd80;
vramData[13'd3893] = 8'd120;
vramData[13'd3894] = 8'd202;
vramData[13'd3895] = 8'd120;
vramData[13'd3896] = 8'd183;
vramData[13'd3897] = 8'd135;
vramData[13'd3898] = 8'd80;
vramData[13'd3899] = 8'd135;
vramData[13'd3900] = 8'd17;
vramData[13'd3901] = 8'd135;
vramData[13'd3902] = 8'd31;
vramData[13'd3903] = 8'd120;
vramData[13'd3904] = 8'd17;
vramData[13'd3905] = 8'd135;
vramData[13'd3906] = 8'd31;
vramData[13'd3907] = 8'd120;
vramData[13'd3908] = 8'd17;
vramData[13'd3909] = 8'd120;
vramData[13'd3910] = 8'd214;
vramData[13'd3911] = 8'd120;
vramData[13'd3912] = 8'd30;
vramData[13'd3913] = 8'd135;
vramData[13'd3914] = 8'd16;
vramData[13'd3915] = 8'd120;
vramData[13'd3916] = 8'd210;
vramData[13'd3917] = 8'd120;
vramData[13'd3918] = 8'd148;
vramData[13'd3919] = 8'd135;
vramData[13'd3920] = 8'd16;
vramData[13'd3921] = 8'd135;
vramData[13'd3922] = 8'd90;
vramData[13'd3923] = 8'd135;
vramData[13'd3924] = 8'd166;
vramData[13'd3925] = 8'd135;
vramData[13'd3926] = 8'd202;
vramData[13'd3927] = 8'd135;
vramData[13'd3928] = 8'd31;
vramData[13'd3929] = 8'd135;
vramData[13'd3930] = 8'd202;
vramData[13'd3931] = 8'd120;
vramData[13'd3932] = 8'd16;
vramData[13'd3933] = 8'd120;
vramData[13'd3934] = 8'd202;
vramData[13'd3935] = 8'd120;
vramData[13'd3936] = 8'd202;
vramData[13'd3937] = 8'd120;
vramData[13'd3938] = 8'd75;
vramData[13'd3939] = 8'd120;
vramData[13'd3940] = 8'd31;
vramData[13'd3941] = 8'd120;
vramData[13'd3942] = 8'd16;
vramData[13'd3943] = 8'd120;
vramData[13'd3944] = 8'd145;
vramData[13'd3945] = 8'd120;
vramData[13'd3946] = 8'd52;
vramData[13'd3947] = 8'd120;
vramData[13'd3948] = 8'd30;
vramData[13'd3949] = 8'd120;
vramData[13'd3950] = 8'd17;
vramData[13'd3951] = 8'd120;
vramData[13'd3952] = 8'd198;
vramData[13'd3953] = 8'd120;
vramData[13'd3954] = 8'd145;
vramData[13'd3955] = 8'd120;
vramData[13'd3956] = 8'd164;
vramData[13'd3957] = 8'd120;
vramData[13'd3958] = 8'd83;
vramData[13'd3959] = 8'd120;
vramData[13'd3960] = 8'd83;
vramData[13'd3961] = 8'd135;
vramData[13'd3962] = 8'd30;
vramData[13'd3963] = 8'd135;
vramData[13'd3964] = 8'd37;
vramData[13'd3965] = 8'd135;
vramData[13'd3966] = 8'd62;
vramData[13'd3967] = 8'd135;
vramData[13'd3968] = 8'd61;
vramData[13'd3969] = 8'd135;
vramData[13'd3970] = 8'd94;
vramData[13'd3971] = 8'd55;
vramData[13'd3972] = 8'd46;
vramData[13'd3973] = 8'd87;
vramData[13'd3974] = 8'd214;
vramData[13'd3975] = 8'd87;
vramData[13'd3976] = 8'd28;
vramData[13'd3977] = 8'd87;
vramData[13'd3978] = 8'd0;
vramData[13'd3979] = 8'd231;
vramData[13'd3980] = 8'd252;
vramData[13'd3981] = 8'd247;
vramData[13'd3982] = 8'd183;
vramData[13'd3983] = 8'd55;
vramData[13'd3984] = 8'd255;
vramData[13'd3985] = 8'd39;
vramData[13'd3986] = 8'd198;
vramData[13'd3987] = 8'd55;
vramData[13'd3988] = 8'd202;
vramData[13'd3989] = 8'd56;
vramData[13'd3990] = 8'd223;
vramData[13'd3991] = 8'd48;
vramData[13'd3992] = 8'd223;
vramData[13'd3993] = 8'd48;
vramData[13'd3994] = 8'd223;
vramData[13'd3995] = 8'd48;
vramData[13'd3996] = 8'd223;
vramData[13'd3997] = 8'd48;
vramData[13'd3998] = 8'd220;
vramData[13'd3999] = 8'd131;
vramData[13'd4000] = 8'd210;
vramData[13'd4001] = 8'd152;
vramData[13'd4002] = 8'd164;
vramData[13'd4003] = 8'd152;
vramData[13'd4004] = 8'd210;
vramData[13'd4005] = 8'd152;
vramData[13'd4006] = 8'd210;
vramData[13'd4007] = 8'd152;
vramData[13'd4008] = 8'd145;
vramData[13'd4009] = 8'd152;
vramData[13'd4010] = 8'd145;
vramData[13'd4011] = 8'd152;
vramData[13'd4012] = 8'd48;
vramData[13'd4013] = 8'd152;
vramData[13'd4014] = 8'd148;
vramData[13'd4015] = 8'd152;
vramData[13'd4016] = 8'd202;
vramData[13'd4017] = 8'd152;
vramData[13'd4018] = 8'd164;
vramData[13'd4019] = 8'd152;
vramData[13'd4020] = 8'd210;
vramData[13'd4021] = 8'd152;
vramData[13'd4022] = 8'd181;
vramData[13'd4023] = 8'd152;
vramData[13'd4024] = 8'd198;
vramData[13'd4025] = 8'd120;
vramData[13'd4026] = 8'd210;
vramData[13'd4027] = 8'd120;
vramData[13'd4028] = 8'd16;
vramData[13'd4029] = 8'd152;
vramData[13'd4030] = 8'd202;
vramData[13'd4031] = 8'd152;
vramData[13'd4032] = 8'd164;
vramData[13'd4033] = 8'd152;
vramData[13'd4034] = 8'd50;
vramData[13'd4035] = 8'd120;
vramData[13'd4036] = 8'd190;
vramData[13'd4037] = 8'd8;
vramData[13'd4038] = 8'd139;
vramData[13'd4039] = 8'd120;
vramData[13'd4040] = 8'd92;
vramData[13'd4041] = 8'd120;
vramData[13'd4042] = 8'd198;
vramData[13'd4043] = 8'd120;
vramData[13'd4044] = 8'd135;
vramData[13'd4045] = 8'd120;
vramData[13'd4046] = 8'd200;
vramData[13'd4047] = 8'd120;
vramData[13'd4048] = 8'd172;
vramData[13'd4049] = 8'd120;
vramData[13'd4050] = 8'd31;
vramData[13'd4051] = 8'd120;
vramData[13'd4052] = 8'd16;
vramData[13'd4053] = 8'd120;
vramData[13'd4054] = 8'd183;
vramData[13'd4055] = 8'd120;
vramData[13'd4056] = 8'd183;
vramData[13'd4057] = 8'd120;
vramData[13'd4058] = 8'd164;
vramData[13'd4059] = 8'd8;
vramData[13'd4060] = 8'd16;
vramData[13'd4061] = 8'd8;
vramData[13'd4062] = 8'd70;
vramData[13'd4063] = 8'd120;
vramData[13'd4064] = 8'd200;
vramData[13'd4065] = 8'd120;
vramData[13'd4066] = 8'd155;
vramData[13'd4067] = 8'd120;
vramData[13'd4068] = 8'd202;
vramData[13'd4069] = 8'd120;
vramData[13'd4070] = 8'd228;
vramData[13'd4071] = 8'd135;
vramData[13'd4072] = 8'd210;
vramData[13'd4073] = 8'd135;
vramData[13'd4074] = 8'd37;
vramData[13'd4075] = 8'd135;
vramData[13'd4076] = 8'd183;
vramData[13'd4077] = 8'd135;
vramData[13'd4078] = 8'd202;
vramData[13'd4079] = 8'd135;
vramData[13'd4080] = 8'd230;
vramData[13'd4081] = 8'd120;
vramData[13'd4082] = 8'd16;
vramData[13'd4083] = 8'd135;
vramData[13'd4084] = 8'd50;
vramData[13'd4085] = 8'd135;
vramData[13'd4086] = 8'd135;
vramData[13'd4087] = 8'd135;
vramData[13'd4088] = 8'd85;
vramData[13'd4089] = 8'd135;
vramData[13'd4090] = 8'd17;
vramData[13'd4091] = 8'd120;
vramData[13'd4092] = 8'd156;
vramData[13'd4093] = 8'd120;
vramData[13'd4094] = 8'd90;
vramData[13'd4095] = 8'd120;
vramData[13'd4096] = 8'd125;
vramData[13'd4097] = 8'd120;
vramData[13'd4098] = 8'd44;
vramData[13'd4099] = 8'd120;
vramData[13'd4100] = 8'd92;
vramData[13'd4101] = 8'd120;
vramData[13'd4102] = 8'd183;
vramData[13'd4103] = 8'd120;
vramData[13'd4104] = 8'd30;
vramData[13'd4105] = 8'd120;
vramData[13'd4106] = 8'd80;
vramData[13'd4107] = 8'd120;
vramData[13'd4108] = 8'd16;
vramData[13'd4109] = 8'd120;
vramData[13'd4110] = 8'd30;
vramData[13'd4111] = 8'd120;
vramData[13'd4112] = 8'd80;
vramData[13'd4113] = 8'd135;
vramData[13'd4114] = 8'd183;
vramData[13'd4115] = 8'd120;
vramData[13'd4116] = 8'd31;
vramData[13'd4117] = 8'd120;
vramData[13'd4118] = 8'd164;
vramData[13'd4119] = 8'd120;
vramData[13'd4120] = 8'd37;
vramData[13'd4121] = 8'd120;
vramData[13'd4122] = 8'd83;
vramData[13'd4123] = 8'd135;
vramData[13'd4124] = 8'd104;
vramData[13'd4125] = 8'd135;
vramData[13'd4126] = 8'd114;
vramData[13'd4127] = 8'd135;
vramData[13'd4128] = 8'd95;
vramData[13'd4129] = 8'd135;
vramData[13'd4130] = 8'd218;
vramData[13'd4131] = 8'd135;
vramData[13'd4132] = 8'd70;
vramData[13'd4133] = 8'd135;
vramData[13'd4134] = 8'd228;
vramData[13'd4135] = 8'd135;
vramData[13'd4136] = 8'd96;
vramData[13'd4137] = 8'd87;
vramData[13'd4138] = 8'd218;
vramData[13'd4139] = 8'd55;
vramData[13'd4140] = 8'd210;
vramData[13'd4141] = 8'd135;
vramData[13'd4142] = 8'd16;
vramData[13'd4143] = 8'd135;
vramData[13'd4144] = 8'd0;
vramData[13'd4145] = 8'd167;
vramData[13'd4146] = 8'd198;
vramData[13'd4147] = 8'd135;
vramData[13'd4148] = 8'd198;
vramData[13'd4149] = 8'd8;
vramData[13'd4150] = 8'd210;
vramData[13'd4151] = 8'd128;
vramData[13'd4152] = 8'd210;
vramData[13'd4153] = 8'd16;
vramData[13'd4154] = 8'd210;
vramData[13'd4155] = 8'd16;
vramData[13'd4156] = 8'd210;
vramData[13'd4157] = 8'd16;
vramData[13'd4158] = 8'd210;
vramData[13'd4159] = 8'd16;
vramData[13'd4160] = 8'd202;
vramData[13'd4161] = 8'd152;
vramData[13'd4162] = 8'd164;
vramData[13'd4163] = 8'd152;
vramData[13'd4164] = 8'd202;
vramData[13'd4165] = 8'd152;
vramData[13'd4166] = 8'd16;
vramData[13'd4167] = 8'd152;
vramData[13'd4168] = 8'd202;
vramData[13'd4169] = 8'd152;
vramData[13'd4170] = 8'd83;
vramData[13'd4171] = 8'd152;
vramData[13'd4172] = 8'd16;
vramData[13'd4173] = 8'd152;
vramData[13'd4174] = 8'd202;
vramData[13'd4175] = 8'd152;
vramData[13'd4176] = 8'd210;
vramData[13'd4177] = 8'd152;
vramData[13'd4178] = 8'd210;
vramData[13'd4179] = 8'd120;
vramData[13'd4180] = 8'd16;
vramData[13'd4181] = 8'd120;
vramData[13'd4182] = 8'd80;
vramData[13'd4183] = 8'd120;
vramData[13'd4184] = 8'd202;
vramData[13'd4185] = 8'd120;
vramData[13'd4186] = 8'd202;
vramData[13'd4187] = 8'd120;
vramData[13'd4188] = 8'd164;
vramData[13'd4189] = 8'd152;
vramData[13'd4190] = 8'd16;
vramData[13'd4191] = 8'd152;
vramData[13'd4192] = 8'd195;
vramData[13'd4193] = 8'd8;
vramData[13'd4194] = 8'd166;
vramData[13'd4195] = 8'd152;
vramData[13'd4196] = 8'd200;
vramData[13'd4197] = 8'd120;
vramData[13'd4198] = 8'd85;
vramData[13'd4199] = 8'd120;
vramData[13'd4200] = 8'd173;
vramData[13'd4201] = 8'd120;
vramData[13'd4202] = 8'd37;
vramData[13'd4203] = 8'd120;
vramData[13'd4204] = 8'd251;
vramData[13'd4205] = 8'd120;
vramData[13'd4206] = 8'd31;
vramData[13'd4207] = 8'd120;
vramData[13'd4208] = 8'd236;
vramData[13'd4209] = 8'd120;
vramData[13'd4210] = 8'd17;
vramData[13'd4211] = 8'd120;
vramData[13'd4212] = 8'd86;
vramData[13'd4213] = 8'd8;
vramData[13'd4214] = 8'd239;
vramData[13'd4215] = 8'd8;
vramData[13'd4216] = 8'd94;
vramData[13'd4217] = 8'd120;
vramData[13'd4218] = 8'd31;
vramData[13'd4219] = 8'd120;
vramData[13'd4220] = 8'd101;
vramData[13'd4221] = 8'd120;
vramData[13'd4222] = 8'd17;
vramData[13'd4223] = 8'd120;
vramData[13'd4224] = 8'd16;
vramData[13'd4225] = 8'd120;
vramData[13'd4226] = 8'd16;
vramData[13'd4227] = 8'd120;
vramData[13'd4228] = 8'd28;
vramData[13'd4229] = 8'd120;
vramData[13'd4230] = 8'd17;
vramData[13'd4231] = 8'd120;
vramData[13'd4232] = 8'd228;
vramData[13'd4233] = 8'd120;
vramData[13'd4234] = 8'd214;
vramData[13'd4235] = 8'd120;
vramData[13'd4236] = 8'd17;
vramData[13'd4237] = 8'd135;
vramData[13'd4238] = 8'd76;
vramData[13'd4239] = 8'd135;
vramData[13'd4240] = 8'd197;
vramData[13'd4241] = 8'd135;
vramData[13'd4242] = 8'd202;
vramData[13'd4243] = 8'd120;
vramData[13'd4244] = 8'd202;
vramData[13'd4245] = 8'd120;
vramData[13'd4246] = 8'd155;
vramData[13'd4247] = 8'd120;
vramData[13'd4248] = 8'd164;
vramData[13'd4249] = 8'd120;
vramData[13'd4250] = 8'd18;
vramData[13'd4251] = 8'd120;
vramData[13'd4252] = 8'd16;
vramData[13'd4253] = 8'd120;
vramData[13'd4254] = 8'd141;
vramData[13'd4255] = 8'd120;
vramData[13'd4256] = 8'd171;
vramData[13'd4257] = 8'd120;
vramData[13'd4258] = 8'd41;
vramData[13'd4259] = 8'd120;
vramData[13'd4260] = 8'd213;
vramData[13'd4261] = 8'd120;
vramData[13'd4262] = 8'd135;
vramData[13'd4263] = 8'd120;
vramData[13'd4264] = 8'd200;
vramData[13'd4265] = 8'd120;
vramData[13'd4266] = 8'd18;
vramData[13'd4267] = 8'd120;
vramData[13'd4268] = 8'd208;
vramData[13'd4269] = 8'd120;
vramData[13'd4270] = 8'd148;
vramData[13'd4271] = 8'd120;
vramData[13'd4272] = 8'd31;
vramData[13'd4273] = 8'd120;
vramData[13'd4274] = 8'd172;
vramData[13'd4275] = 8'd135;
vramData[13'd4276] = 8'd48;
vramData[13'd4277] = 8'd135;
vramData[13'd4278] = 8'd149;
vramData[13'd4279] = 8'd120;
vramData[13'd4280] = 8'd16;
vramData[13'd4281] = 8'd135;
vramData[13'd4282] = 8'd207;
vramData[13'd4283] = 8'd135;
vramData[13'd4284] = 8'd17;
vramData[13'd4285] = 8'd135;
vramData[13'd4286] = 8'd37;
vramData[13'd4287] = 8'd135;
vramData[13'd4288] = 8'd210;
vramData[13'd4289] = 8'd135;
vramData[13'd4290] = 8'd145;
vramData[13'd4291] = 8'd135;
vramData[13'd4292] = 8'd16;
vramData[13'd4293] = 8'd135;
vramData[13'd4294] = 8'd94;
vramData[13'd4295] = 8'd135;
vramData[13'd4296] = 8'd214;
vramData[13'd4297] = 8'd135;
vramData[13'd4298] = 8'd16;
vramData[13'd4299] = 8'd135;
vramData[13'd4300] = 8'd83;
vramData[13'd4301] = 8'd135;
vramData[13'd4302] = 8'd80;
vramData[13'd4303] = 8'd135;
vramData[13'd4304] = 8'd163;
vramData[13'd4305] = 8'd119;
vramData[13'd4306] = 8'd198;
vramData[13'd4307] = 8'd135;
vramData[13'd4308] = 8'd230;
vramData[13'd4309] = 8'd152;
vramData[13'd4310] = 8'd183;
vramData[13'd4311] = 8'd152;
vramData[13'd4312] = 8'd202;
vramData[13'd4313] = 8'd8;
vramData[13'd4314] = 8'd202;
vramData[13'd4315] = 8'd8;
vramData[13'd4316] = 8'd202;
vramData[13'd4317] = 8'd8;
vramData[13'd4318] = 8'd202;
vramData[13'd4319] = 8'd8;
vramData[13'd4320] = 8'd210;
vramData[13'd4321] = 8'd152;
vramData[13'd4322] = 8'd210;
vramData[13'd4323] = 8'd152;
vramData[13'd4324] = 8'd210;
vramData[13'd4325] = 8'd152;
vramData[13'd4326] = 8'd210;
vramData[13'd4327] = 8'd152;
vramData[13'd4328] = 8'd210;
vramData[13'd4329] = 8'd152;
vramData[13'd4330] = 8'd210;
vramData[13'd4331] = 8'd152;
vramData[13'd4332] = 8'd210;
vramData[13'd4333] = 8'd152;
vramData[13'd4334] = 8'd202;
vramData[13'd4335] = 8'd152;
vramData[13'd4336] = 8'd202;
vramData[13'd4337] = 8'd152;
vramData[13'd4338] = 8'd183;
vramData[13'd4339] = 8'd8;
vramData[13'd4340] = 8'd202;
vramData[13'd4341] = 8'd152;
vramData[13'd4342] = 8'd202;
vramData[13'd4343] = 8'd152;
vramData[13'd4344] = 8'd202;
vramData[13'd4345] = 8'd152;
vramData[13'd4346] = 8'd248;
vramData[13'd4347] = 8'd152;
vramData[13'd4348] = 8'd252;
vramData[13'd4349] = 8'd152;
vramData[13'd4350] = 8'd200;
vramData[13'd4351] = 8'd152;
vramData[13'd4352] = 8'd210;
vramData[13'd4353] = 8'd152;
vramData[13'd4354] = 8'd230;
vramData[13'd4355] = 8'd152;
vramData[13'd4356] = 8'd249;
vramData[13'd4357] = 8'd8;
vramData[13'd4358] = 8'd218;
vramData[13'd4359] = 8'd8;
vramData[13'd4360] = 8'd84;
vramData[13'd4361] = 8'd152;
vramData[13'd4362] = 8'd252;
vramData[13'd4363] = 8'd152;
vramData[13'd4364] = 8'd75;
vramData[13'd4365] = 8'd120;
vramData[13'd4366] = 8'd110;
vramData[13'd4367] = 8'd152;
vramData[13'd4368] = 8'd48;
vramData[13'd4369] = 8'd152;
vramData[13'd4370] = 8'd212;
vramData[13'd4371] = 8'd8;
vramData[13'd4372] = 8'd169;
vramData[13'd4373] = 8'd8;
vramData[13'd4374] = 8'd202;
vramData[13'd4375] = 8'd152;
vramData[13'd4376] = 8'd28;
vramData[13'd4377] = 8'd120;
vramData[13'd4378] = 8'd74;
vramData[13'd4379] = 8'd120;
vramData[13'd4380] = 8'd16;
vramData[13'd4381] = 8'd120;
vramData[13'd4382] = 8'd166;
vramData[13'd4383] = 8'd8;
vramData[13'd4384] = 8'd155;
vramData[13'd4385] = 8'd8;
vramData[13'd4386] = 8'd198;
vramData[13'd4387] = 8'd152;
vramData[13'd4388] = 8'd84;
vramData[13'd4389] = 8'd120;
vramData[13'd4390] = 8'd16;
vramData[13'd4391] = 8'd135;
vramData[13'd4392] = 8'd200;
vramData[13'd4393] = 8'd135;
vramData[13'd4394] = 8'd210;
vramData[13'd4395] = 8'd135;
vramData[13'd4396] = 8'd202;
vramData[13'd4397] = 8'd120;
vramData[13'd4398] = 8'd202;
vramData[13'd4399] = 8'd120;
vramData[13'd4400] = 8'd16;
vramData[13'd4401] = 8'd120;
vramData[13'd4402] = 8'd202;
vramData[13'd4403] = 8'd120;
vramData[13'd4404] = 8'd230;
vramData[13'd4405] = 8'd120;
vramData[13'd4406] = 8'd214;
vramData[13'd4407] = 8'd120;
vramData[13'd4408] = 8'd197;
vramData[13'd4409] = 8'd120;
vramData[13'd4410] = 8'd159;
vramData[13'd4411] = 8'd120;
vramData[13'd4412] = 8'd17;
vramData[13'd4413] = 8'd120;
vramData[13'd4414] = 8'd202;
vramData[13'd4415] = 8'd152;
vramData[13'd4416] = 8'd126;
vramData[13'd4417] = 8'd120;
vramData[13'd4418] = 8'd200;
vramData[13'd4419] = 8'd120;
vramData[13'd4420] = 8'd16;
vramData[13'd4421] = 8'd120;
vramData[13'd4422] = 8'd183;
vramData[13'd4423] = 8'd120;
vramData[13'd4424] = 8'd171;
vramData[13'd4425] = 8'd120;
vramData[13'd4426] = 8'd92;
vramData[13'd4427] = 8'd120;
vramData[13'd4428] = 8'd95;
vramData[13'd4429] = 8'd120;
vramData[13'd4430] = 8'd92;
vramData[13'd4431] = 8'd120;
vramData[13'd4432] = 8'd18;
vramData[13'd4433] = 8'd120;
vramData[13'd4434] = 8'd162;
vramData[13'd4435] = 8'd120;
vramData[13'd4436] = 8'd37;
vramData[13'd4437] = 8'd135;
vramData[13'd4438] = 8'd48;
vramData[13'd4439] = 8'd135;
vramData[13'd4440] = 8'd129;
vramData[13'd4441] = 8'd135;
vramData[13'd4442] = 8'd171;
vramData[13'd4443] = 8'd135;
vramData[13'd4444] = 8'd148;
vramData[13'd4445] = 8'd135;
vramData[13'd4446] = 8'd83;
vramData[13'd4447] = 8'd135;
vramData[13'd4448] = 8'd16;
vramData[13'd4449] = 8'd135;
vramData[13'd4450] = 8'd248;
vramData[13'd4451] = 8'd135;
vramData[13'd4452] = 8'd214;
vramData[13'd4453] = 8'd135;
vramData[13'd4454] = 8'd80;
vramData[13'd4455] = 8'd120;
vramData[13'd4456] = 8'd198;
vramData[13'd4457] = 8'd120;
vramData[13'd4458] = 8'd210;
vramData[13'd4459] = 8'd120;
vramData[13'd4460] = 8'd67;
vramData[13'd4461] = 8'd135;
vramData[13'd4462] = 8'd248;
vramData[13'd4463] = 8'd135;
vramData[13'd4464] = 8'd183;
vramData[13'd4465] = 8'd119;
vramData[13'd4466] = 8'd198;
vramData[13'd4467] = 8'd135;
vramData[13'd4468] = 8'd210;
vramData[13'd4469] = 8'd152;
vramData[13'd4470] = 8'd210;
vramData[13'd4471] = 8'd152;
vramData[13'd4472] = 8'd210;
vramData[13'd4473] = 8'd152;
vramData[13'd4474] = 8'd210;
vramData[13'd4475] = 8'd152;
vramData[13'd4476] = 8'd210;
vramData[13'd4477] = 8'd24;
vramData[13'd4478] = 8'd31;
vramData[13'd4479] = 8'd152;
vramData[13'd4480] = 8'd210;
vramData[13'd4481] = 8'd152;
vramData[13'd4482] = 8'd164;
vramData[13'd4483] = 8'd152;
vramData[13'd4484] = 8'd209;
vramData[13'd4485] = 8'd152;
vramData[13'd4486] = 8'd164;
vramData[13'd4487] = 8'd152;
vramData[13'd4488] = 8'd83;
vramData[13'd4489] = 8'd152;
vramData[13'd4490] = 8'd181;
vramData[13'd4491] = 8'd152;
vramData[13'd4492] = 8'd80;
vramData[13'd4493] = 8'd152;
vramData[13'd4494] = 8'd210;
vramData[13'd4495] = 8'd8;
vramData[13'd4496] = 8'd210;
vramData[13'd4497] = 8'd8;
vramData[13'd4498] = 8'd183;
vramData[13'd4499] = 8'd8;
vramData[13'd4500] = 8'd90;
vramData[13'd4501] = 8'd8;
vramData[13'd4502] = 8'd17;
vramData[13'd4503] = 8'd152;
vramData[13'd4504] = 8'd248;
vramData[13'd4505] = 8'd152;
vramData[13'd4506] = 8'd209;
vramData[13'd4507] = 8'd8;
vramData[13'd4508] = 8'd210;
vramData[13'd4509] = 8'd8;
vramData[13'd4510] = 8'd183;
vramData[13'd4511] = 8'd8;
vramData[13'd4512] = 8'd212;
vramData[13'd4513] = 8'd152;
vramData[13'd4514] = 8'd31;
vramData[13'd4515] = 8'd152;
vramData[13'd4516] = 8'd210;
vramData[13'd4517] = 8'd152;
vramData[13'd4518] = 8'd210;
vramData[13'd4519] = 8'd152;
vramData[13'd4520] = 8'd135;
vramData[13'd4521] = 8'd152;
vramData[13'd4522] = 8'd166;
vramData[13'd4523] = 8'd8;
vramData[13'd4524] = 8'd95;
vramData[13'd4525] = 8'd120;
vramData[13'd4526] = 8'd250;
vramData[13'd4527] = 8'd8;
vramData[13'd4528] = 8'd124;
vramData[13'd4529] = 8'd152;
vramData[13'd4530] = 8'd95;
vramData[13'd4531] = 8'd152;
vramData[13'd4532] = 8'd210;
vramData[13'd4533] = 8'd152;
vramData[13'd4534] = 8'd106;
vramData[13'd4535] = 8'd120;
vramData[13'd4536] = 8'd214;
vramData[13'd4537] = 8'd120;
vramData[13'd4538] = 8'd210;
vramData[13'd4539] = 8'd120;
vramData[13'd4540] = 8'd210;
vramData[13'd4541] = 8'd120;
vramData[13'd4542] = 8'd202;
vramData[13'd4543] = 8'd135;
vramData[13'd4544] = 8'd16;
vramData[13'd4545] = 8'd135;
vramData[13'd4546] = 8'd109;
vramData[13'd4547] = 8'd120;
vramData[13'd4548] = 8'd31;
vramData[13'd4549] = 8'd120;
vramData[13'd4550] = 8'd171;
vramData[13'd4551] = 8'd120;
vramData[13'd4552] = 8'd83;
vramData[13'd4553] = 8'd120;
vramData[13'd4554] = 8'd230;
vramData[13'd4555] = 8'd120;
vramData[13'd4556] = 8'd90;
vramData[13'd4557] = 8'd120;
vramData[13'd4558] = 8'd16;
vramData[13'd4559] = 8'd120;
vramData[13'd4560] = 8'd159;
vramData[13'd4561] = 8'd120;
vramData[13'd4562] = 8'd17;
vramData[13'd4563] = 8'd120;
vramData[13'd4564] = 8'd202;
vramData[13'd4565] = 8'd120;
vramData[13'd4566] = 8'd16;
vramData[13'd4567] = 8'd120;
vramData[13'd4568] = 8'd166;
vramData[13'd4569] = 8'd120;
vramData[13'd4570] = 8'd16;
vramData[13'd4571] = 8'd152;
vramData[13'd4572] = 8'd28;
vramData[13'd4573] = 8'd152;
vramData[13'd4574] = 8'd28;
vramData[13'd4575] = 8'd8;
vramData[13'd4576] = 8'd209;
vramData[13'd4577] = 8'd136;
vramData[13'd4578] = 8'd39;
vramData[13'd4579] = 8'd152;
vramData[13'd4580] = 8'd80;
vramData[13'd4581] = 8'd152;
vramData[13'd4582] = 8'd200;
vramData[13'd4583] = 8'd120;
vramData[13'd4584] = 8'd31;
vramData[13'd4585] = 8'd120;
vramData[13'd4586] = 8'd17;
vramData[13'd4587] = 8'd120;
vramData[13'd4588] = 8'd30;
vramData[13'd4589] = 8'd120;
vramData[13'd4590] = 8'd17;
vramData[13'd4591] = 8'd120;
vramData[13'd4592] = 8'd135;
vramData[13'd4593] = 8'd135;
vramData[13'd4594] = 8'd90;
vramData[13'd4595] = 8'd135;
vramData[13'd4596] = 8'd83;
vramData[13'd4597] = 8'd135;
vramData[13'd4598] = 8'd30;
vramData[13'd4599] = 8'd135;
vramData[13'd4600] = 8'd202;
vramData[13'd4601] = 8'd120;
vramData[13'd4602] = 8'd210;
vramData[13'd4603] = 8'd120;
vramData[13'd4604] = 8'd80;
vramData[13'd4605] = 8'd135;
vramData[13'd4606] = 8'd172;
vramData[13'd4607] = 8'd135;
vramData[13'd4608] = 8'd210;
vramData[13'd4609] = 8'd135;
vramData[13'd4610] = 8'd80;
vramData[13'd4611] = 8'd120;
vramData[13'd4612] = 8'd75;
vramData[13'd4613] = 8'd120;
vramData[13'd4614] = 8'd202;
vramData[13'd4615] = 8'd120;
vramData[13'd4616] = 8'd90;
vramData[13'd4617] = 8'd120;
vramData[13'd4618] = 8'd135;
vramData[13'd4619] = 8'd135;
vramData[13'd4620] = 8'd202;
vramData[13'd4621] = 8'd135;
vramData[13'd4622] = 8'd76;
vramData[13'd4623] = 8'd135;
vramData[13'd4624] = 8'd183;
vramData[13'd4625] = 8'd55;
vramData[13'd4626] = 8'd198;
vramData[13'd4627] = 8'd135;
vramData[13'd4628] = 8'd145;
vramData[13'd4629] = 8'd152;
vramData[13'd4630] = 8'd210;
vramData[13'd4631] = 8'd152;
vramData[13'd4632] = 8'd210;
vramData[13'd4633] = 8'd152;
vramData[13'd4634] = 8'd202;
vramData[13'd4635] = 8'd152;
vramData[13'd4636] = 8'd210;
vramData[13'd4637] = 8'd152;
vramData[13'd4638] = 8'd16;
vramData[13'd4639] = 8'd152;
vramData[13'd4640] = 8'd202;
vramData[13'd4641] = 8'd152;
vramData[13'd4642] = 8'd210;
vramData[13'd4643] = 8'd152;
vramData[13'd4644] = 8'd210;
vramData[13'd4645] = 8'd152;
vramData[13'd4646] = 8'd16;
vramData[13'd4647] = 8'd152;
vramData[13'd4648] = 8'd202;
vramData[13'd4649] = 8'd152;
vramData[13'd4650] = 8'd202;
vramData[13'd4651] = 8'd152;
vramData[13'd4652] = 8'd30;
vramData[13'd4653] = 8'd24;
vramData[13'd4654] = 8'd202;
vramData[13'd4655] = 8'd8;
vramData[13'd4656] = 8'd80;
vramData[13'd4657] = 8'd8;
vramData[13'd4658] = 8'd80;
vramData[13'd4659] = 8'd8;
vramData[13'd4660] = 8'd183;
vramData[13'd4661] = 8'd24;
vramData[13'd4662] = 8'd214;
vramData[13'd4663] = 8'd8;
vramData[13'd4664] = 8'd210;
vramData[13'd4665] = 8'd8;
vramData[13'd4666] = 8'd210;
vramData[13'd4667] = 8'd8;
vramData[13'd4668] = 8'd202;
vramData[13'd4669] = 8'd8;
vramData[13'd4670] = 8'd210;
vramData[13'd4671] = 8'd8;
vramData[13'd4672] = 8'd83;
vramData[13'd4673] = 8'd8;
vramData[13'd4674] = 8'd183;
vramData[13'd4675] = 8'd8;
vramData[13'd4676] = 8'd210;
vramData[13'd4677] = 8'd8;
vramData[13'd4678] = 8'd230;
vramData[13'd4679] = 8'd8;
vramData[13'd4680] = 8'd207;
vramData[13'd4681] = 8'd120;
vramData[13'd4682] = 8'd16;
vramData[13'd4683] = 8'd120;
vramData[13'd4684] = 8'd85;
vramData[13'd4685] = 8'd120;
vramData[13'd4686] = 8'd230;
vramData[13'd4687] = 8'd120;
vramData[13'd4688] = 8'd16;
vramData[13'd4689] = 8'd120;
vramData[13'd4690] = 8'd80;
vramData[13'd4691] = 8'd120;
vramData[13'd4692] = 8'd80;
vramData[13'd4693] = 8'd120;
vramData[13'd4694] = 8'd202;
vramData[13'd4695] = 8'd120;
vramData[13'd4696] = 8'd31;
vramData[13'd4697] = 8'd120;
vramData[13'd4698] = 8'd202;
vramData[13'd4699] = 8'd120;
vramData[13'd4700] = 8'd80;
vramData[13'd4701] = 8'd120;
vramData[13'd4702] = 8'd70;
vramData[13'd4703] = 8'd120;
vramData[13'd4704] = 8'd202;
vramData[13'd4705] = 8'd120;
vramData[13'd4706] = 8'd80;
vramData[13'd4707] = 8'd120;
vramData[13'd4708] = 8'd208;
vramData[13'd4709] = 8'd120;
vramData[13'd4710] = 8'd183;
vramData[13'd4711] = 8'd8;
vramData[13'd4712] = 8'd83;
vramData[13'd4713] = 8'd120;
vramData[13'd4714] = 8'd179;
vramData[13'd4715] = 8'd8;
vramData[13'd4716] = 8'd95;
vramData[13'd4717] = 8'd8;
vramData[13'd4718] = 8'd34;
vramData[13'd4719] = 8'd120;
vramData[13'd4720] = 8'd252;
vramData[13'd4721] = 8'd120;
vramData[13'd4722] = 8'd16;
vramData[13'd4723] = 8'd120;
vramData[13'd4724] = 8'd252;
vramData[13'd4725] = 8'd152;
vramData[13'd4726] = 8'd94;
vramData[13'd4727] = 8'd152;
vramData[13'd4728] = 8'd191;
vramData[13'd4729] = 8'd152;
vramData[13'd4730] = 8'd166;
vramData[13'd4731] = 8'd152;
vramData[13'd4732] = 8'd34;
vramData[13'd4733] = 8'd152;
vramData[13'd4734] = 8'd94;
vramData[13'd4735] = 8'd152;
vramData[13'd4736] = 8'd248;
vramData[13'd4737] = 8'd152;
vramData[13'd4738] = 8'd17;
vramData[13'd4739] = 8'd120;
vramData[13'd4740] = 8'd31;
vramData[13'd4741] = 8'd152;
vramData[13'd4742] = 8'd7;
vramData[13'd4743] = 8'd120;
vramData[13'd4744] = 8'd16;
vramData[13'd4745] = 8'd152;
vramData[13'd4746] = 8'd95;
vramData[13'd4747] = 8'd120;
vramData[13'd4748] = 8'd202;
vramData[13'd4749] = 8'd120;
vramData[13'd4750] = 8'd30;
vramData[13'd4751] = 8'd120;
vramData[13'd4752] = 8'd17;
vramData[13'd4753] = 8'd120;
vramData[13'd4754] = 8'd198;
vramData[13'd4755] = 8'd120;
vramData[13'd4756] = 8'd135;
vramData[13'd4757] = 8'd120;
vramData[13'd4758] = 8'd16;
vramData[13'd4759] = 8'd135;
vramData[13'd4760] = 8'd210;
vramData[13'd4761] = 8'd135;
vramData[13'd4762] = 8'd80;
vramData[13'd4763] = 8'd120;
vramData[13'd4764] = 8'd188;
vramData[13'd4765] = 8'd120;
vramData[13'd4766] = 8'd252;
vramData[13'd4767] = 8'd120;
vramData[13'd4768] = 8'd76;
vramData[13'd4769] = 8'd152;
vramData[13'd4770] = 8'd31;
vramData[13'd4771] = 8'd120;
vramData[13'd4772] = 8'd164;
vramData[13'd4773] = 8'd152;
vramData[13'd4774] = 8'd30;
vramData[13'd4775] = 8'd120;
vramData[13'd4776] = 8'd202;
vramData[13'd4777] = 8'd120;
vramData[13'd4778] = 8'd80;
vramData[13'd4779] = 8'd120;
vramData[13'd4780] = 8'd252;
vramData[13'd4781] = 8'd120;
vramData[13'd4782] = 8'd16;
vramData[13'd4783] = 8'd135;
vramData[13'd4784] = 8'd210;
vramData[13'd4785] = 8'd135;
vramData[13'd4786] = 8'd51;
vramData[13'd4787] = 8'd135;
vramData[13'd4788] = 8'd164;
vramData[13'd4789] = 8'd152;
vramData[13'd4790] = 8'd202;
vramData[13'd4791] = 8'd152;
vramData[13'd4792] = 8'd210;
vramData[13'd4793] = 8'd152;
vramData[13'd4794] = 8'd210;
vramData[13'd4795] = 8'd152;
vramData[13'd4796] = 8'd164;
vramData[13'd4797] = 8'd152;
vramData[13'd4798] = 8'd210;
vramData[13'd4799] = 8'd152;

