// Testbench for hcount module

// Assume that #1 advances time by 10ns.
// The test bench will use #1 to mean one clock cycle,
// which would be a 100 MHz clock, even though in reality
// the dot clock is 25.175 MHz.
`timescale 10ns/1ns

// John Winans's tutorials (https://github.com/johnwinans/Verilog-Examples)
// recommend this
`default_nettype none

module hcount_tb();

  // The testbench just needs to control -RST and CLK
  reg nrst, clk;

  // Outputs generated by the hcount module
  wire hCountEnd, hBeginPulse, hEndPulse, hVisEnd, hBeginActive, hEndActive;

  // instantiate hcount module
  hcount hcount_instance( .nrst( nrst ),
                          .clk( clk ),
                          .hCountEnd( hCountEnd ),
                          .hBeginPulse( hBeginPulse ),
                          .hEndPulse( hEndPulse ),
                          .hVisEnd( hVisEnd ),
                          .hBeginActive( hBeginActive ),
                          .hEndActive( hEndActive ) );

  initial begin
    nrst = 0;
    clk = 0;
  end

endmodule
